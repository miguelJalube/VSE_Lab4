-------------------------------------------------------------------------------
-- HEIG-VD, Haute Ecole d'Ingenierie et de Gestion du canton de Vaud
-- Institut REDS, Reconfigurable & Embedded Digital Systems
--
-- Fichier      : avalon_computer.vhd
--
-- Description  : Sequential calculator on an avalon MM slave
--
-- Auteur       : L. Fournier
-- Date         : 19.08.2022
-- Version      : 1.0
--
-- Utilisé dans : Laboratoire de VSE
--
--| Modifications |------------------------------------------------------------
-- Version   Auteur      Date               Description
-- 1.0       LFR         see header         First version.
-- 1.1       LFR         13.10.2022         Correct behavior readdatavalid
-------------------------------------------------------------------------------

--| Library |------------------------------------------------------------------
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
-------------------------------------------------------------------------------

--| Entity |-------------------------------------------------------------------
entity avalon_computer is
    generic (
        N        : integer range 0 to 32 := 3;
        ADDRSIZE : integer range 3 to 16 := 3;
        DATASIZE : integer range 1 to 16 := 16;
        ERRNO    : integer range 0 to 10  := 0
    );
    port (
        clk_i           : in  std_logic;
        rst_i           : in  std_logic;
        address_i       : in  std_logic_vector(ADDRSIZE-1 downto 0);
        byteenable_i    : in  std_logic_vector(1 downto 0);
        read_i          : in  std_logic;
        write_i         : in  std_logic;
        waitrequest_o   : out std_logic;
        readdatavalid_o : out std_logic;
        readdata_o      : out std_logic_vector(15 downto 0);
        writedata_i     : in  std_logic_vector(15 downto 0)
    );
end avalon_computer;
-------------------------------------------------------------------------------

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1_1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
PdDOWTu+Lr8ci8Pg9vMNnqbfh71HZpxyEVGdDRGlFj85JKZxM5e17IgNtRm53Te3
fF9vO2repyPcTpx/gkRYe+NoMqDg/d336iGN6bQyXCLyxUXY0yoNuJuMRhW+AMFV
aRuw2hf4KCUL733WChALkj35huoUH6Do+O9kcNn1MwMHpsW/zwX0X1GWmjEKJBa7
fe5ZwmSkw3dAb+1/P+PS+ZBLyBTRIW3ehJmsIpTaeQ+wvAvU9YQW4ItdpsehI9vg
KCOgIUHzM+sG5NjZxrYsN7Hc4Z0VemvP8MmEkrtkXhefXm4NNKyM22LVRVxWn/Z2
oc5qLgZPe9YHRa2HL2cgRA==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 20480 )
`protect data_block
PxdqtquOgNnlQRJASvv3FZODH3qqa9+Md9xNdGUNpYe03yMWVm+7bKwrBNmc5Un8
fSI2gWPtAIrOS3k4vGFVdXC8OnrS3pbkLM15fM0HIdK4YUS8qFPw0+lpDNGqQEh3
Z/zPobt3hXR+dbBRmNIQRcS/iL2WQmbhkudhZNER/iB/2RFHW3EnTWJXTJmFJqnY
cIkhdxsg0SURVoXeDUEu0LMOcPHgXv+RWmSmyOTN/w9md2ezSvwdVOdSphqDKsyc
eWDPZgLoY69NGX1Zjw23aNLPWVuHpea4XbQQe18tbAGqbFJQfuRYnCBsq5MjXKqn
4z1t1g8W7pj0OVWwTKNppdw14tuC9vVgVEegyBtKgfjTSAWjPZb4ze7H0Upf/NRn
QbCKeQCP9/2NzC8aqwo5Ey2AyKfnOCius6EI5UMFzRxnimYQ0ujuI989ex8q0K1j
GxZH0yA5L+PhnGRYFm5JIG8S6vMXmMfIEv1F2vYMz0WDiOaYSeOjYW0KI88YwPFQ
iMeFI+PxXEvelsMRRzf3kxrQ0/I5zZ4ll3ZvpxAU13U3NFWjLt4RjT42T+/cTWe3
fKs8FWKJOyho6h2WToh7VRE1YBw993MNWgLQKVw71s9HOEwssrRuSy7uh+6f3pUl
iBf9x6JqRXOvMt/ye4Cq4YKigYeMmy7tWVLYB8xrhTL3bjzroDgtf6oUYBIYsiEg
4EeNlNcJUYWWD2unhseqdDaDs66qCsE+5wohBFwQdI6njo2/yu+QAXFXsK5oBlpL
tn0DE/8C1rVoAIT72X9S53cC/82NxmC5lp2w/vkVfxIj5Aa5eZn6J3I7XdG0ulte
/vVfKoag4gudpF4bAcCegMSWiww6ZTsq4swtXxlXB/WKOBUDBLuq5+6QNkJkTTRO
Ajqo5atj3+amMv2K6OJMR9E0QbQ1eemUNsc3fFRyE1AlE7ASZ97S2XbZI9Yjj3IZ
aOlsZnTyyb+HHJqUVbFpcAukyDFxmNnTvC1BhjEM9TfO28dFcIFATxlMtjbmxZOS
3MPJT2B+45asTlOv2wxgehZDwK8W5Xd6nNg3SAZcmwyRfoFmh8astQFIS0qDH2O8
aRgDqRaVoVv4JheUDGeEtAnDnr88JZaxhQhj6wmQv6C7XaHhQA3iHMu8a5f0dBk+
Esa0D3qJFZibgMCdiWmNgSx3ixUBNTO/9t82g+mbZExe3TtVoYH8TFJ2/8evRhWv
dyU5n3LvMruk7SXWRB2rXjGTiPyiSj6Ty9f9hmNkDCEsdmIhHqOWsRVwSjLtRXP1
1qnPKRnuFg1tqMFsgV6ckZTqoRf8CGb7rhliGFQ1NydNOYGjAteLRcSNTH3h08CU
cui1xaGrI5Th6gFgtn969mvXOdz+1er575bD71sEtuIFpI5XypXMrqvpgSTNYch8
WIo+83WsRU80gzA+zAOUBbkUeE3gmtU8p6rR9t5ls4thYnArHsIvhR4UxixDl0I4
ekTRyzZF6ddeGr/kvYarEIHNNhUDQURj/jvAosBwMEE/dEOJch+s4vh/bpO8nK6O
T+ThInNqHxCt12bnBBgzEueeJ7x4uon8tXgeT1tE79B3R9xTEc60Uc8NVUuXWDfg
JkSycpvt3CMcDQetTOlEB27sU918VftGVuKyxMr1FEabO/x7uHTUl18upoNNT/PU
TKFiQscb7FH9YyLgyMr4xZipcuQ4IO39Hnc3bus1/yvf2yeaJC7//aXzis1AJkpu
jeeVKuZQ3Thc/kdRMBMzo1m5z7mSbttscG6VKFYV2KdukAd2vQ+U2C6pxsml2FFy
IVeDp2QhZMlCFhVNm6RtdRbrgh3UA2IgjhQ2iaG93LcOv6ntlMWi16w/nI1Q6i6G
xtRdTUJiWHTZC3hBq3CyshzeK7LcoRBIoCa9GwCY5HC327VrTt3rKgm8r/crjiUF
FVuOwoEaPF9PiLzvfKK+LOUu9ZiCKoMavKxL1y03Rb+WSFwKCL52fq2T2sDC7jjg
lnu9iFYAr7JpK9aDPT5NpySfZHFhOwoW+nuq3Xr9TZqETAyMOtroro55gc1DeOh/
OFcI8ygytivkRV0QbROJfM3gPXfTyItVOWWJc0c4LicneqCDTpPjjUmSkjOQEmeE
QB3x6yUk75xBTF21ezLcbeffnH0A40uCf0RAk2wW0/RnIVBIV64oJh1M08ErZLYO
eKQGHfZ3Ys4ICNCfppB74R/aNxtcDw7B9v92xvb1Hvby04n9WKdOgwi6qHBLDxu1
7bDJ8qvNnXFxVJHSZImIKaOx92jscETSzcADPvoBISci4qM4OGj/3WGFE+fE5uKG
AvbBpBwNN+gODshnkI60JemFCVFSpM7Nm6pDpeEOjMsSqHNpsQepWFxrRVzdQVkj
96q9eXvlzBYmW8vQ9hxgUuz9+/lJT6VFR5eJZpW5u70nZ4NqEXuAnTOUZdSpbb9q
5cVWc13F+T/CCF2CsI2ys7sJaTUl/Y1D653XT7fju3dn+32gC57RCdM/nIG0Jzza
gAZaHJj63sLnoDqfsR3L4t3bVqzh1S1xr8W1SFD2I9hX01bgnXx1rr+OGd66EPJU
guBrMoyWNIcfnll2/HauSyhgbZOpgR0f5K4aUxlnPnE4Un/1xWwvtU3TI/5qQHSR
o0NoFSPK+AZYOII0+9om8kSMy9vIOUVsxxUjlqJIttpHtNoXi3y+t9dyPH+kDtRw
zVaR2n4vHMfjhJ4s3Gt9QsQxYp7GILAq7qKNXPK0KsyBOVFgyeoxbOo4qLzywxvy
Io0j8ej3cmfcDneC1sJ305/OTLjn/PSOJACnZr6Mlni09QnC9u9C43QWw9vJP5JC
zPn+acIjLtiqX5MTgr491LiQIWKcL5vYecTAHf9mSsrQM5WCsYC7f/F7X8KAkIYv
cfaCDW/GwWFbM+qxcu2c350p11h1hPMYx/6F4PbMTNd61DxQCxG5/aBPUm+WJaCs
V9XGPcgv9XvWPXMdlHBeGClyFCHqioLKdPOkokAS7J/7JdOiF1rXPcRyjXTzVgNW
lmjAGgOtPRN6GcsW2B93Kdp5FNX/reuariPWt8V1PUy2ux7+nPZQjWQfsSs55MZd
MUUUBhWfIu4ug2WqiMOkFx9wswcDYzZyzPLet5cOkuZHq9ZeqLxwF3Fztdk0hCGE
y7p8i+0O4m8fsWJ1L2vd6p1zO/9G15rw0O0Roz9SP2eREVyYp4/D2xayekdCFXhV
BIsYuzbhHdiUSmZJCjfINQMUKHhz+R7ioT56JQ635qe/XXgQBH9WhxdpMcoWhqOD
kma63uUudJ/pO/ZIgLBKaKCx2KZpEEmFSTYsnRG8HJjWn3x7FwvkLZp807DHXJQP
NOfOtcRh2Qj8QhuxhBqcFL73UvtBp9VK1XRNVL60a2Rpm3HLjUIy2zfY5WC4OIhU
E+y25xmEc53LJCux+U5bOCkMIhL00heMAzDd2qDg/yLwlOsZcvfP1WqYSoLpD4W/
DQMNXN4RKjCwEIhvFtpeMtbqxpy/Rlm8+6ieIAAQ8VP6+Xzg9CTnOWTrgZtvaDVe
dLOKz32tjTJj4SBHxVHaew2ZlMrj8Uk7+qm9s3SyIW8MVUiX5JBOMz563nHIiuS+
zAn4DB9+ZmX8Aejja3ZjueMc903kPNxuuUTPket3NVLdh014KIw2IrWuxbotfMy4
Hq/MtgDTKy1y9eUMZsPi19S7sdY01P+020LjXQDM8Ysgpt0Wa3sRyxDwhs/lGTtI
rXvltpUxyGz9oygUGabAqByOMP6/Vt2l8hPBXu6JG4Nhbsp1qUEw8CJ7uiZJsJVk
bsjW+NzsrDNyuG53lg+KLmOWpOQAXd9+1PtkC9yXRSWZc/Rm1gATwv8v34MfbsMq
+1bMzolHNgyLQOisyEUdk+9mUlkxhw136BwjE8dWClseaB8KLc03+WmQZjhvIYxQ
YRblajIjGXEZydM62MBlC4ImGObGSaIAumTFCHgRYZWTNTprkhhI0rl5Whxak3kr
duaEX3OUY9CY+P4JwUwRZqkjPnrDbQrNPDT7ohj92JrgZUl1ltA8gMuJE/sjDM0K
NFoQNje3i6/PWV/HihKrbS+uoZfMvO4BQobmSVFDpx0YON70L0rNdJar7kI5oY9F
kJKEii2rJE1XEDZ264PwJqKYAutrON/ZKGQWGCYPdisFHHS/NaXw3CcfujNU1K3u
qacOI+EdLeOxJvyR7nFIflIovdVYXQRwPc+GOF5gDRUNz+AQpWYjKZPnYpFgxreD
1sdJnKNzGmudFMUUdWIEEr/jeTVK9f8qfumCqBmpOzss8j6AF2BIkHnU+YGIZcp9
7IW9scQt1/NQ4ftSAgBsZ/IIuGGL6Hwc2+RAmwofHXYxd06QPvrSc/STwaYOtOnW
cWsLoq9GdrdYplTPquNjVZ2wYalg5gqCBlAN22dl+Xj95Xpn0TZHiRsPFGfSVgqt
cmeuPzNI/Be/fwV89POHFnrp225mLRcbGb1lLPlc+Fk+JKkgUL3aEgPg6+woqKu1
CPw2je4rqAYlozcQlZ2fDnxuA5qwh9VOD3NudviNO9RkVXK6SgBE3kS2QYx0/pmr
11MGUszG0wE1o5VhNkCYtqz1kSoRmmjLHY4o+D060kHn6kOaSAcz6XHR0BO1KlE5
9xxacYSyOm4HQXGesZPeey0PPGwnbplFJX0yPdnZLpu2I2cj/Nx9JRYK0/PLCpxp
9OHHD6xc2ZJ9ZbI/bKS24UJCbgRTVa5DTYCOBQaxV84hd6uu2IbhZWmHrsO73SR7
ewGwnGGywQC290i6T/FhyPdxlIup0FY01LMTfcA81CTEANjKREiQzPf7Ds13btdF
UN+ji9QFKMxgmNMKlP3MAGH5fDVj3hJUT91dMmAsZjRo+KLb6wVC86qnXDoulo/g
zjBiwuqklbAQnV63Zmy/yqkGm5/xKu/5eTVRvmZaUZ3pEDCi1GyyAS/VnrJQFu/0
5wWuyX7bzUISdQ8ji41J7ZqqcQYtX0RfX6NJVkAxYuUtDajKeOEgxWrFnvm6KugH
KLKVnLf6pAxRK4AsUcwD4/CZcl3TtyrSLvomyvT7GAfiTEmjw0jNhRQCjOPS+xQR
grgOzmDvm7nPw14C+AsnlXEjX7/BYB3dxO7LfhbXRi4zfoVgq5c+905JSifWk9ZA
VDPKV5q03v4koY5cxTxZgYK/9i5plGa8WqhPrWUW9Y9vO+EgdTc4yZUd+t28lVzM
KqH8YcmwUljM5XFo5rPlcTT7UeprjHBOtwiv/vqe39MzfeS9lUR81SpHaGQJnol+
kKpbAOEtAS+GbMAoZzEdD78jB6pL6vIyTfqEgwchDOl0fHVjZlBEwmJ83wuQQdtg
ApghPsIi3Iq+RsrjVQ49mMYpg2/iOCXCb1TnTKVOOdSDAqp3hOC4XtZgu8CenuJ3
m9aOGT9OjGmyIygpDOzsI2jL4ltA13elAlc8Ne1ccdsmjNxcjKsLBwhoBuh8yVxZ
+HqDeiwPQtYqBiOc9LFg6wNKk+iMC4slBovxX/onHedvooCKeo6yfWWa0ox8Xo/N
7fS757FrESHNQWZqociDMJoP/F8jJL1WZsQBQ6xQ8aIVr+sR0gD0vdfsDONiHHOt
t3YZdJ737wQdq/XCML0OWKcaZzccU0U1ouVw6PQTEobQc8GQk9EtGAl2t0ah4gpQ
XV0RwDYXMr5H0zddYjHtYSptznsfqQSACdrBI3fbxGwGLY4G2B6EiqHRKXtL+gaj
1SBkBtgURmuyCeFGeP0HpVR5IkO4eVbZ2E5u/UjbSk7ArZ656z2D8qYBzPGaWKvY
DOtXIxUldAjgakHMH5Lsxkr9YxEloM7oeeFlOczrbLFWEoB8qIWN7XwAymt4SIjK
QQEvrdsifRl+3KTYUd+ERlOpLKdMb/TuhbtkZgIIr9FJ/Grkt4dWrxdLSanQqeyQ
XuIkAWUPm61CzdSwsrmMfJ34c3ecRogkVZh0JCm27+zv5+nNcuxI+MiiHkCtEGaD
kjwLBTWqHouzKbQ26UDLWSSPSP9rHPCSQFt6zrRkiVRtnc5pOnYbdvwa3lFMb5wW
UqTOhl0BJxSwmm5n2esPEghhhUoYAq5ajWaEiIMrkoRlWuEXku0WCJxHVwh7/qF8
E5M5J/Njk2Ucs+dIysKH9TbnBfxeGyFHgd1CZVJglsrCtUqfWSZYwszpqSFB/2u1
2DHWgX1fk2ErweU+LVv9Sr87yVjWrtRmQ+vU/eOb0mWzZgM3GOjgO/PgwPgPTdMm
FgK134bYlFoQNFKdOt1vFZhguQXtIJ93JkRY/nL8r8LJcuMVz/ZdZILi2qH4/l6m
BHKHxXQ1Edsd5ZykzYdwc1YZqp5ntT7xf9FuP78NUfdd37+7pzP6ONngJxVkwlju
Z7G3IZxI9O9edhgc5rC8dSEems8H9hzkNL7tefj5Rf52xzoVPv+29Cjv3ud7iyBi
+Sty/kdJo3ShMkgmhF+3Fy2GhvEMFLQ0lY+DkhQxg6CqqxeT+ZNWdhyytLGF/fDL
MRYWIhw7s832ZUd+i75ZDaDE2hkuap7+vq+O+grUh6m69WBgQJ7hg2XrvbUzHqNw
hHQSbAN1lzMy3cjcfq6Uukv3Gx0xOqfgVvrR/ARTTNKqS56vYWQ1DfGuQe/dM0dy
ivBJ+3LjhAaZNMebJlPw+v6LkLgExu6EeBaGVuFevnipeY1CuFmb/UuW+UjEfgPi
CVcNGEdhHhZZWmgQn0d5DyigrAYlhsqDdgszXLhrwljLDR3rkfE77Dt1VpoQHPNp
sjWPYB5hyneL65gdpbJAMzZu2eJhunmb6Ldmozw8a1p8/h9W9uaainRwyvfS5Wvl
h21J8NypH4yf3wfcCIamwIOgflEzT33yuFrZIY4whU2j6e0Pm359RB3rlmIuZJZ9
9PeHue+li/HUUccDpoVP0Qk7SsOVT9JT4TVPqlimzGEZqX9NLFO+6XC6fFRCp0kg
a2fUEDG4+u5lztq+YkCBXAsl/zD3ePD6nDpslhOcHeQ/19oIyIAsBoganOj5QFFl
K+DedF7VUDpbwDD5OUnQGNwxLlYU9mjTLDADUhAfwwXGVPIddrtOruRJpY12yrye
AE+JQ30b77TzoQ5zJEXLwqzDMVvtLvWijEwhZjm3+erF9hxl1K/T7zYa8FEu1SKd
OLZXM+nZGbIhPiDYvG3UpuXYQw+V6BPY4PZ30cr4C0VQDxWVsHFpskczV92s82sI
bsHaG4f4M4MHnoVtXcE8gXo6tnkMIFlWpKsvgvEfax38gqqDafpiaQGe+8AXo5m7
IfS2ZHBCqKJF0aQ6w2sfwBYJO4FCtH3eKbMd9Pkwt5AjDFjc5SRSherKkx29d3Rs
fSMQrmOgP8LGwlqpqPmb5jvMIygIbgi3gHvaaTcXtnYwIm1a2CfEm5OEVvsnyJkJ
6PBra5SfEjRUcGQ8ko7cickeF5VaWLaV6BrCBajzvJeYDFADnGZyqR8G2MQELhbk
/9lgQ3GsF4HFz6VhAf38BXtYlnEeaGZa+UOZinVUPlACskNxzkbeiA+P1TrbR1XD
8q7kVamASghnu+CnOKA34p6LtO0EYcbA09yGb7A8DGzeU12iAWnGrjDGUrC2qtbr
htig54CQVK1L1pKallhtWSB8cgSMzh59hrcLz500JgLbuDm8bixR4nCJ/2vtcLV9
oJPcyZK5RXM/m4pzl48G1JeQHTVb8x8EH+im1tjn5ZSxnDtsKwNB5z2hOrYX3Phc
ZJx35+bVERCw9V0BtgOAyt2td94GlGrnvRD/tzTUeEfE4IkZd+chz+Y+VGN74iYR
ESyVOv5butUZgsYXj24J5hJMdRXV0wrfTDx33UmlduIlNokW/QDHvORnwYqpxW24
/pQ8nhVGvfFprqHcFTMGYYoz3BVvzZJUO0gZeLhjSqu0MX+mfheMYC/TEKZVbMUd
g7YadfjDm8fzHpsTFhNR+Oj/nVVqOD/XGyfYM00KGhgz0jMoEqN4+wwAj20z6aDs
ZZo0vMY9+JBNqm6I+VPHV6H1p53xP6DK23aVGjOepioo70gf2MOYpBv9QaZJm/zZ
BL58zKc8ZftScWwMg4ZTOW3BL6kYwxPxfe6m4SqaWyjW3VXGe0Bi5hsFSnir0GQy
N205XGCo87LzokwzJ0lteXb6UR2Gkhd88L9ezlZqgAx6oKrQHXlqYgDzX/4f75JQ
vDYRsWgIjVt7CV5gEMb3eYi6e/h7cQlCmk6odiA+dNViF/HWJjA5Jm/Au0lIzMwQ
gWtIzXSNBfySzZIWgPCLRacF8yRVo2om+lzZw1D/XIQx9U+gY1TLbkg4TW3iu71h
ebmq+94xJjvcD7kcnceEabw+HbnqYK0Lk50VMwWH2iWzWAmiuepaYQBmY9215vqj
3ZYxhbHZUlqAkFZdjg+fAu9VWNoftjilwuNOygCGulOEyw05dQWQ/yW1/flyCzFG
hjd9S0MSe52Dq7eQMJhhtwxRsmIlwKTSJsnuE1BXl19nfje/TRAEteoqmebyDpAo
zCyP3FAfTXPcXB5uMOgeuUMByqEt/+sIIfdn33fvSPxAAqxpH0/wxB9aBzotJvnl
I7xxOcJBhfJJ/xSlOfXA85JRBjvtpqOzzkn+/3X+aKwG/Gyp2+/ZhN3cTDriPhKR
rjv23+Ib1aGfpddJJgJBElil5LioJYwf1ShrIlU6YxZKImnpPBHSBSh+d3AMA0bG
M+eUsss6kRugOFpqZsIwjyNRhgIyZ2EZNcbUkOOnkHEQciwt9/DeL87+pqUwUwuv
yahYc0QafWawCdUqnX1ya886NmSotK4JC4HNXPzy//3OGJaaSd9R2pKKMl36FvgA
7B0BKIm+GAH7fxRWxtKKV/cEfcxb5qRm3/bollP90VkyTmgF8I2CHI67eIIevaNk
Yt5wOkfbZaMfAZuUJFP1d55aH3n5g8ypmTIxlpcJoB/MFVsV4Be3fO9V28CjPCXh
6ggEoC5aF2nk6hrz8RamOrWa1lBONJJkt9cWBvHtV5AZptyRz4WYbnEW2ryWZwlB
3I3T3MJtmHw/tU7HOCYb0YB9DV4xhsHXO3towkvRbLyhmBZK+v/DR0ajn1dTW06x
P+eqZitIp4rNa4c+Yq87zBJzOEEnfFryFV8lcRzPDtHd1zFQcQPH/nQ+tpGCIF2n
EjmNy+TTL0Yvov+JArFkhfQQ+jEW5aYExe5DDdlO/tKeup4CF2bTCns9+4cfl2Fn
rlVzzF/h7vVu6yX9xUMaFIr2IWWfK6ipMAGkR4IbsWPh48IDimDvqPK9qqzh6Gm1
EG7QUzZXOlAD2gXT1H5IRoJWvCzVjHhqYlc77dgu7jbRAehXUgYBUIbf8034PIzZ
Cp8N0lyserBXdUJgvSjZyIEziAjUzPY9RQCPBJZ0T5eYKpiu+GbHoRJHGjncVsDi
C4qM/HDU2ej2UxXaz7T8BJEXxMZrzjJTab65PsYl52G4RaZwXvM27w0Mug1y5wI8
xsrbwK6ey9mOxTXCP0aAs3BQYfPT1VSFfClR6PvKt4LA40kxYr4H8hefnP6Yu/We
4R8lyL1qCSzXy0C/85rUq0UEmttHsY6Ch6+3nExYBCvCJmad0De1OlI0sIB86+cm
emrnqNqZbthjPCvHKRkDApM/ZnxHWTSR0x08hf8RajaD9L3v47MZe78ORO7NdcBM
WiWna6WzfHLNr7g1znhH995l6MxOPZVRh6DIABbiF+FzKXRRNL7gjGnYPjqO7Dq+
Nmy1nFLxW2nH5/cCAcmK8GOjMCKAjMd3RNqEcCMbiUajfaDU5uBM3ZUh+bV6ZV3Y
yL2noU4nb9vTO6PeGQPyCK8FK0V+Gue40+PewhBJofXpeM2naat21AAPTEcS6aP5
jY/zkDgoG4ksbpadz1q8J4A5BoZHCrHnUhbbe1V+mcdJTYFIcI8FQjbXDQtXLgZI
jSeVubRf/i/hNV1zOWFTZFobXO7+JBrlLSJTL1jSsPntxaF17AWP21MyXRuqJ4C2
v4lwFiCyhQLUSyBX3Uxt0yUFAcR0iMDK0p6gmujJP1SEAsAy3segEG1QufdeGwko
1iffBGPhltYAvUYxqLoYWzlVWM05lZVGih+hai5FaWznpmw7CFHz3/bHTB8G4PEU
0yxD2SiaRss1JarDWgTjJJ6wp3g89T+LPzRyGpFhpq/C0OVhNt6sNJ/VUlFFu7ct
JPL6EGC0l55kQPMRuUaziFWhQQ76NB+WVAbxoVEt7TOFES27iv1wBd8T/EdLmLzP
0WiOhBGyS0pdCCuFt36ETqQcQWxgnLTup0vOHGf84pTwNL5lnHZC7a+aV3qs0vUt
NsKS8rsQ50fnfIbUtg6hdrZEZI9cr/BW4T0v8TJIWgsey1Dr7rnGdtqlBum5515T
QKl9Ie2kZJKy7eXhbZtWDv5/XlqDnNRfByMK6UgQRIPgFKqUphuJdutElC2q9xJZ
ruwPsqwacV/5AR6N1YzahoMX2Q876jk21nyOvmQXyKybIpELu6atBLiVkIRanBTX
tgrlpjvyN0exCxkpyw5hmkRyJnAfUlJvO2LulWqodGGKtfeBQZUVmDh9VFIJ3z0Q
/pJ8bhWa+s4FEpacIhcmcli7rXCrvZWhsgnPRb1CN3UUhhs7gUWnT8UoRUEFnNmV
sNiBMgBfuipFiYK6w8XZglLg8gfIgAc/qkDj/x64KlV7GnCySlSTDBc3WgxWTNUT
HT3Qh5jBD9xBPy4GTuO5p3fIsVg4pLzwLF4HEyRg3hHWrQ9nTsm/Zk/FDZQbYBC/
pje9ITkfkl/kuA8Qbbs6zjZLBRlq5rh8Ne5FvhyaDSfeaevn5uHfUOpG4nnFI5Zw
YNQVn5S7kaZ4XzAXmDj0Xvfmp4ayTq5SZf7i39WxHm9wKK59nBQQmRU+2yszdnoK
jT76ghPh+ANfxCX1SoQq0aBUtOIkFr7KhAALwL+APlfJKd4L9wPMWTXLua6lve+U
0mS0s//GzM2ki0AaZLVZo3HBXfVMO9keFD4v6xHStKr833CnvBWm3fv4YhqUDoAt
5wixdcZ86AEEYBpL5Zq3jjr7Met0fwVyvWDXlelw+2E/VNjHibL0yRYGy0gn+cBt
kRYa60vuoq99m0smkS6w7PAgW7UUK/mQPEzsgdu+z8pqXU4qmFPfX7ahjeL2qN0I
VziNEpNv/Zy+GGdK/21RZxEN28EGFw77O7Im/ufeQRpsQT+Elgrjt7MCounGUqk5
UJR1TpLX/hXIf5vSy3TXwFtLHxa0R5Xdl+Lhd75t1ZMFb1YGfm75Jg4ywyqAJ8jh
R4kK1A0CgGh45AUIZfo3GWuAUEmaJI0U1bR2sqNc9p11J8z0U5Ko28zv5FmaiLcr
sSb362ccB4E2VjQvio4QYahncX1TrR0zFgx2+Z+GcWryanqJQsZC50M90a9Ql5nr
BNNa8aRyeG0ZBGyB/cPwJCR5aojT6BCL1VtFJmqTBaaF4nIZMhfFYkLTQgwtXICH
E/PRTFbomaXARa872YOTcUJ7sGVBuFIJU2eFIwxJHZ2eA7u0ytr/OQzggGJRU0Ch
hfRIqcRwPSokSRPnM0nM6gTLlZ94EGFOqZRj93+pP1NLjdtX09btOQ7oJwwCahKT
TS9wayG6LPODAykbKLpft6NCBi/NfrebmdCcPSNKwS5Qd7mf8tQJvwknDQQCAdru
7x/H3arSCt3DWOFUYWqkeL6Vo5QXFvwNiZGxHWgVxxS+BpJPGLh6eYv6hzBzPWEy
m9CN58DbnhTjE7kTCNcNHIQkahejnx4a3EUEtFT9O4vzb0Z04kKcWj0L0snKFb6e
zY1/rZxGEbIOdV+L6FdTzCTRyvvpxkWXNHKvokWA2YuJ9bDzLPxbU4YQ+3x4/9d/
oL/LKxIwYRGWXHRk4R+ZqxQovnQlE8/DjAfMvhwavrohNiia2NJmHn1jRNZF+bHN
WbcYlMi3bEj9OOZSeAJPHMBZHV/SO0YePwZf4zBimf7ea8Ibd+bqxtVoIuOvR+lu
/tkxF3t797eR/xlHcGFci/x4veb9p50GG2K1oR1EfhwgKfD/OZfgWpo+eJBPxh+9
Xu5zDzoF5zcq2Nfdc3u8L3d7FTXLCaXB2rmS5B0dcE9krx9MMEnCveRAQSxnaiDR
oq99aNgO/w2ZAz787XjMHGmqOUBKg0mjEszSB9kFgoeiQNVw2GiYp5mtkMfJVT/L
cu+6KRHlnu65MsJ39LEgG/ImwyinKHnUAIWIrCMPbrJTZcOl96An1sxZLFXAXmil
ksM8yxtAv3zDRVVviKv0tSRykMaU69SitJ9gNa5ghr5J2WJps8szjsRJa9pU+baD
3+wxs0IkHTYIOmk7JOfNm3odHzuaNgHdKremKWnYjby9VCN2cbaA2bLaIWidOU0D
mVhK8vybjtOFa4XQu2US/VlAQ5RItVMIy9qCVff1Fl9pwKdVwt6x6FCNE8/VSmU8
N6J5h1q5ePlNJc+WBlYkfr5w9mgEdEYGtNg6QJqMmVAdi/04QNUvG9HvrQgvctZP
wztb2pN293Kvs2AwBbDAI2kGWugIxjAR1aClsTCh0JUK3/DRqeOs8dAVIhan1qwo
R9WOvhRWoVR5kEm3WojOXAlsSelNV6JfolCLFzH5WwnE1pOrmhwfqrbwEYMybp6y
m9u1HdS32WIdy7Berpr7iO9Ggdlz9B/Qh4LpVDUMl9Ot4BGLK8nXPfJTjlkvwYsm
KX+wc9bmoYp3mG0ljCBpG2EyRzmCwc+ao+63y1xcHeyRjCY4MvIC5uXrYHeGLa9a
xyjSL8ia4h2biUL/U1pEORxcFxzvSQIVw320U1pgcJjbE+6DuZEgchVT33mEgNgw
HAuUCzcz17y+/jxgKgLyUrv3GKRjQI009J1bUf+c8626ZxJGuGneb5TgsbfKEgF4
HGax87sZHA+fzELvGQtKJoM8JTKjMiIZ2wU7aBGIBU3pXESSL5Zgx06LELFCRMKw
C40SAMYqs6Nn0DJeJcGJQucwBXKEIikgWiVtvtMKHlolwb+kEjBIAj5sH02vWBCk
kRJCggIB9DKUMVRj3RcFbcIfxFbS7vun/9/0OPSRUfg0o54v9/J9zftYQvu5F43C
9m/WSUoAqDsWVomv9wIFGVRil/JNQCBNl3MB60DN2xFeH8qpP/8Lz+lFKUoutEOX
4mcBFAhiLQdDYklqJ/4KnVdNY2H/OhMs7zFRGkkqlLAEdjmaDPaT2xgaQUG+9Gse
UJugRJYGgLB1AuoI+uoOPxN1R5JiVNnaBQE9SJUl5h1UxUu9ETl45lb0frM0/F0j
0/4lhEFZDvpRnSwQ2Fu5Xwq47PfEeh0LT75ExqhIkwfYyyfjVgqn77oBTcvYUP5+
b/tjMjqwSAmVcsMAAPBxfkgQ1LrPBzWv0UbwdKAO1VWfzpdTE9jhf1A3MuUDMjlO
+c7gcFuwe3D1g0rmvaQE0knDhloOuq1k10aeRsU7yhVZi0wCO0JyUlDMRLcp6Fqi
EkHaxnzsTxYmjwUOPNdFt14qru/gws1HZIj/+SLaoAjM5IGRkwLiSUSgE5HJLcH7
g3D/8hMfIizXcGEyX7kgQX8Yk2ILff/L5eBFfr+JuxxR/Q8gZ8n1LG0zXaYF6RNy
xabfT5Kk000pvzkwokWADUlqJEksqwimxUJFWsSYmTpn5eg52b10ZE545BjuYney
I0vYs9cppAGWT11Q+QIdAL1p+7P13mW0WocQTKZUDX2SN3zo/vsIss13tIdMK8tV
/HPB9EyhgsdWXf8jDqNcyVibl7gY53uggtCGVXAImCc0KgOL0kKm95elmYcYrT2O
6n4I4PFDMMpx1vHkddzY5gUo/qsj/8c+HihND2RpxyZ+HyeUn0tlMnshmH72T9VY
8PimW0+UhIbYmUabj62byFGqkSVkMBeTqA2oV7Hx/eNqQLNFz7evXxOnkPanNbY8
TR3C93nwdRSATJjFKBvLBCyM5r/Ckc5VDjKl507Nm0713aEy/Vgl0zRwwqargFrt
uIx9OLyW/BQ8hw/p7UcqSU5R1BRFL+m13BdVXOpJT5IanFWQqcNLWblIpM3x1JIa
c8a61YEA1FrvzSYizbxEWDc4SGFjEWO9oU9/CpJ9A66Ha3kFvZTMugXaO8FrZ7ip
l8oM8U5vWXhRajT0Nvce3OGGFmYUJVvRB1MMVR7MOL2nsLan//54w98+XvLwrE10
irAzH4NWCdBHvutR4Q04GZX4fdtBD+VnP/rMwlYeMXAkdh4ic1GHKWkzlLvs89TL
cRW14Mds9K5X4RaJtN+JwTw1QyezolnPR5kxLacMHM0VaDvQmJS6Okxqv6hcmBP0
LSUiw2YO9xWudeScTX5Mkq5vqltPFpczjBoshxCUZdqL7bkUzEFKhoSg6cdYY4CN
SXof0J6nt33IZ7r/V2J+XXvCrOYEhdeQcCazXzvONoPcolODlmVl6Om5toUC+Hyt
Kyl6vGP32BrVfQ45Fr2abN0AXiNZaFSrDV+8c6OzPNNrmjdYZ92fwELkbTvwMY4J
6lq9A/Fcpr3Z94sie7p+rUYo3zSarmw+WA+vf3Na9koNFwiusfQVFhdkc0Ud8toh
58LzI77ydKNmX98gEGD9yDrqcY7QHVs2v8fs9TLarbiwuSSZPDrIE0AN3jmUwguL
QpqoCo7WNANoRWpbVSMcWyvvx2X+5u+pA+60VekNJti5oY96kXZEKfztNade714k
u7Vx8mtgbhtL+A8cZfOpG5Tu7Tw6kImU762NQlub0y+QM7qBfxST6Sj08w8CbsJu
bUZrD2cd+iXFdcM1egUOPRUYMMDNZvK/DF2RrDgooQNtqvIrMRxSJoam7iX2vO+Y
FOB9qhcZo94bpp6imgGgbbVs6+0soYGfjR0SOqfuVlj5PbNV/ryJDdMorIewrQ52
u0UFCZFY9t7GH/yty6XV1fATwm9nabNJLrw6v2m2YKJ9QzcAKjbMnjhGoL+T+Apq
9BXBGJJ6qqSc7NOAQD7AYnBX13k1aG8vfqlA/VdNoDEllpRSpyuMUfjudFUlkQx7
ez1LPW5p4XfUR1KVAIhfQe5HO4+EssZ7/WFuLCwWq5C4he/+sNZhsaJN1ep1Mint
CQQOnRBoSrrIU5DzUM5dNNP4gqSlUxn69Oo0sNn60iLGcNggqySvHnx5lXbS3lQE
3JHLv5QVAlbO6Zxzy8ZZ4oWHydKvN2KP5gAnsTxAPlQsEKBvyg7LGOhJm8Zd6ge/
amN9aM5UBedPavL24Pof75Q67+X+xACyXLWEuQMnZbbZtgNOV3G8H98+fAp+DP3a
71Osy4Z1Veo4G+fE3bOZ3ED4bxi1k87oYVP/4dbs2yrF9UHvwJsoCRlkKXhRbm6i
OF/MGaCM1RMw9RIlP/pka0Cl/wXmWn8PoMblx9mi9m15IC/mWmeLgJwggl1zAnTn
gQXkOsuoXOmPS9L+LXJhL5+I3wVpQK1etJAsf6vN7p9fXoluhX47O9MbT2vTIvp7
VwjhMXnLwOJIulSQDnJfBp2ggsD/vZ2vcTD80ZrRPp6zsc+i2fQtjznjml1cDuN1
SYptRqYYnBNS9Zw9erb/rEKLur8gH2c+710adhpzPOjrpHG6oyl8hVGMOtXL4z7E
W1hIio/v7kFzzk2IhxHR7eXJJusvYOEnAEjbZraedCYCkByegXWE3IPqrT2UIIlK
IcSmgEjhCtfxRC6p2C75BuuaZOkZDCLy6Yh6TcnPGlSZMQsgIGqmSNl4Gbwj0IN9
NqZJXxIljvjRgUbiNOj8It6vk/HpjIk0NxYk2g0pJG9j02H84x4KXHoPv0aIJgiw
t6TsAd9dzOrfO477ajf8FLcgsjFE7ZrUf6h7oNfjsGVWE+4eUBBj/gkr8+ILBQ6O
dXKltOcoHiH4TzGWluilGzM3AWupI4s3I7A8Cw8bVg3V3q5hv8bkjlGIMkxTWK4N
dszygSZvauALrzkkv8JRPrWUlcCl2loHAFcKISmmQgoy0JEIc6VoBh/Uu7Wsh2T9
CPHMko8UbWeVEPDDVAUtblFyVQfUI2RLKPXrOmpCp9kFPwpgjZqV6pemtjSkfGkF
5l5A+8Xz/yLpci1aK6g3dhHHda4haT/82JdTV6HS7lrgV857880waZNo49E7ibRw
Ipmx/C+jh2gpnjddCY6qTkDLpZcvf09FftfsYtmI95P1er0Egthy6uYm7n2ckZrF
iTkiAa57KUGPvMOGQkA8Qx6Qn0SPEiOzkxW4YxmxNalHW6FC+E0NyXE2hfCAcj6j
BNmzCQaSKSmgD1M8iyehykhBot6yixDmclFTXOxbK0ICYoe57PLfKGNgMU+RVDYd
mmxRw4st4DEYvmabsYOe8dbJR94a9oVNcF06MapUvoXoq1gokG6/Z9Y+tRBrjzza
Gdrs5OYwjG94HB40mDfAuUjIFDJNiCvOL+l7XgMeYG4JWWsoQXHoV18YH5ESi0QX
M9A4NHb3QR61YC1odi1/rKN5N9UhorK8awXOW+rXFJkIG6ZPp9Kl1Y3UHgE9m8GF
0XFQDoykDF3YqObJfDFKSLbdFVeZTp3/2gJbeF8Px1gBXqdY++me9xKQ6v4rDzPO
afrAC8lKxZ4XpATmpHujvS2fVhsjWldFMGHFonixl+71KiKRLpoUEsDSlYpEsgsN
nlAJAMrim5Q6wqKMgMc8eoOENUj7/7xuUvrGxXBkmOWl0gJsW6JKM2VboFobrYZq
ktsMJZg724W8Z+4dV6YRlV5ef9Vk6qlbQkHCMnHo+cIWFoOtBUZVrEwqCMtL++QK
gCX2yeMdcnV6cqT7UcNMxZNLbUJFCm3oKfiW3WjLlEpP5YXe5c/Kdfd5VUkftIKC
ggEhTlirdN/YiGfDBkUU60LHsbgNRCOFoQDZd8oCtgfnEmWOD48X8Lt6mbY748as
NWRPI7cOnFaxf7fbFFa/0Dr3uqj4w5WIHCx+WpyINLWb5/yPZhMQogW8BqX6sIHo
YnPT1Ne1P2amHZvANxEtoO+VMbzGPVvtJldKTtBk4tD9cTVXBBZJyv1aZj5Ytqsn
BHrCvOB0wVKKRRbTQN6aKHAyprDubI1EpZACjUat1/0s4LyEGD3UuXmEOYrcSYwg
6JV4Oe6R1/rfIz9rzSbQFuTsQtXIfd9FiW5u54porCUS/4jUCGY2gNWpN/gmFNHZ
Twelnh0XNTmjUsRsgt0toeOsT9l8Roci/2slrR/VMptBYzqXzvmAHiXJbsb132h6
XY2cAkh/O3VHcas1EE2gfZj3PGk/Tj54Anj8hdMIEwPcmsNT6gYdDVQHJzCVsTfI
YYoio6F7JkhycPtc31TwGWBPHajlKW/pNI25ugt0PlXXNt6uN5lQUHQeJsRQouaS
YxeCPDYfEuy/zs8/g9Lp2FvbXgViXtSgu0zVANCrQ+2TSmtHVCNRtRxY9aivRE2L
3CB9r8O5KlCWmTJJk1hPgoS5N08GySrHEqU76k6NnSTyhSMm60wXbt7NLDmebIVC
NCPKMyf4vtJzvqyu+bRsKA7yA5Kz18YugHW9xodK2DNDf8JEcdzSHlGZZY3Gt0fP
cNMwH/4Nugv76emZpW9rNsL7pdy9ZhaHWY/SHUVjdOqx3uflNTz/cWe2zs9K9sXf
T+182Dz0HPKgIX1eJKL+8P9ItyvL3pDCI3iE0FX/Vsd2NIQaV2NgWSGzWSmYA153
uksqYWQzWUCZR5fuMRMyPfCtkvN8mwt8bjKy5RlmYc6yT1d7JrfQp1926Q3aR57D
0n2i1q320C4bePfIh1LxXSbAuvMYLlWOQNv3EEiJ3u3t6UVirjyZJrS33VXjd2lM
ZDWIHG4o2AeaTFSmne8Fy+O1OZfG0mBqpSZjis2eTPnf/vWb+Qc4KzY2KATZsV4w
46NSjaZxZjtsBIjy70H/sN+qvDzPWTO6SynYDYqQespf+lf0T3FmSPq8BmWLxH7K
X/H+/0FM7sNMb32zVrQ8PHL3oxbdWXU4ZlnoRuhIQ2l3IeGdRaizRCWa9whVBoK8
n3OyH0wK0yPj7CK2TNcpPMDqMhc9WlUK33xq7S0KfiyE4qH5T/YOXwQ6kbYRIflH
RTWz9I5jn6rUtH0BTMtVb5B3Nvn03ftIWU36vPKVY5RffoLYnnMHzFB2TnOAsBzW
ikwZJ8B2HQHTBHHOx81cYsVk4jzFNySDzkm+wbqqKFwf81imuMmZIn47j7xhaKQB
JOCUKo6dqj07wJL5APMDVkVl0kgRTPJTdgYy0J7GgktOXFWKUzAejH+UAtzyv72u
+OEx05sWkjIn2f1vk3Ucz6UQMUad/vvKIPZTrx+v0pnrUzfyOADvofdMIaOEf3N4
VZVypcsBWYt+mkOACxOg7rr8sjXvKLqECb6nB39aJeh5RDtbbb+M1f1GO8urhEU5
dZtcIc6+LdpID/wZy8CGy5w/RXMhzttlb/FCL+5338N/rJJMhxXijvGudCjCmZxi
Ow+sV4uLOtY/fSIbKEZLEx4Jjn+R7z3KYaHArXmCTh+DQquJOI7OaR25E+USNSy4
HL2Zm+zQyQzMnj+1MLrtilieSwnDaXVWfMcLhewV+aGlUes+7NOOV8IPZCfC9pU3
V2gVfeNkNX8WoMiaJkstrpW83NJNxU2LR8D7iM4x9jZBWrqXi5B0keIu/HDkS/87
6QzU6MYnkiaBqcUP2u+wX4TdQCUsEvAwSB6WrLBrazN2v8LZgcIyyQrK8NYm/N1v
/a08vzbhv5U9I9aUAj25J1P6qOyzXJs0l+U12zAkRYnDpDNNeckpgWPR+NhTSDxf
g8RaFKGj5lFV0M1yc/crf1/rj6Au7mPtC0pVeLtRFsxwtvRUoq0Ztr2Hpoe+ORVE
VRAKcHAAQ4LFdXHi2NOF76RVvDgurPzXMOBy/aCYbW99nJeg9T8YK96ixbUbX9ni
kirFoC6AhZ5wX+EPMOX8xN5oWbT4mIVdeCdXVx7JfhR/CzLyWhk5mRV3RUGWRBFS
fm9LC9apS2OLKSG13sP3Gczr4sYfRkNmqD8O773Efie9NMqN4Z0P7is6F4uNvj6r
9B06bJyZ5izzRqC1c/1p/ZV1razJV20B9mz6hmRz+o5fgZbgxLuEDAabhOhjvcUZ
LPPlQ08VUudxiMtk3A9zshQtTa40tsMj9uX41ycrmAc1yU7XZMEEcoNRuM564eR7
x8lTM3fb3I+GFFj3MJ6ceNj8cuA8x4acXRWntIdXewLsQldvxunV/NO+Wrlk/bcb
wDZM49e51LXOCaTR/wA0XHX1+FlyYj2wiYrh7HVj0PQKY3sDmDnTtUlZrAT8KLq9
/LK7lzqKG5nsNzIprFQFxcI1gI1IlxNzgyAqubbrwePMQxOb+9Zut7xwviVFcP94
uurIHFdzqHc7sAhSVfOnY/Jg6z2k7CPTcrOXVdUsp8/lPQ64sSmVLH5KPYotJZTb
goO6fmEh7e2FQ4yLjAINjSzJgR0IP4XxPGyxy07EdSjogSRNtX5Qmp+xjP8zJ7S5
bgVh9ng2ICD6ETBOjrulen7XE69DLGi6Osmh8Dn6a1rgvdyRUoCuVR/CAT30ssN4
OJsnf+Z36ZYVrjgeWRTqKU+iId4xjX3oOOqdH//jSVD7zATeGpx7HCaBuUFaTNkJ
x+ttlsBiP3BHopiYJT91A/hu1eUIsdqDGK/tOEhqnemGEpv0SowTfPkJM6SmAXwi
F9tOCo+N8OCOS5pGDzX6arb0ykmiJPSEL7wspCHYxFc65GUYm2HVfjCsxyWw70xT
w2C2CE6qJlemtkIMp+3PEbiaG7DQDKDsHqW3yzq4KB79HEdIjUNnaljmFCbxqxW1
vTiwMy6BOw2poncz2AFcdJJLtyiNasoIl0utseGEziFso5aKgumrOTqbq69uWLIV
gedYVNK7ccJfH0KSg56+wdHG3J66pcuNGY7/MfbYIBkG303ovBJuOCenPRvl6upl
ihFmsTr0VU4qRDRPWd6jxYNcm4XaCk9Muac29mSxAJEqwrEUlXiMArtiFnlNTEbQ
/65Q9qY1WXRZrhyo3u0q7sACzerXZOVb23ee/SMXpcJVcp/nTa4VE2uIBbBSKbxj
hNCehJohVS/rPhh/Urd21bHj3k0CfKauOr5hv4kmZrap18XoPQVgqLjxmUowAboW
O5UbsY4IjrbJWk2xTL5KZanXrGoCGb1aJ3sVFNORyDxluxG54wOHzfQ/wVEuC+qd
UAmA1+ossvLXDXopccfD1gfKcxrhfd+xm83xvggRAWyZ2fZZt4qnNrWD3zzFr+XK
VQfmGWbgCNcMS8fsTvA8vZ+RvCCoUD91uIKsp1Was60FvZyjOQA3orArohTVjzel
/KIh9kxRfOl+lmCYTlrKb33pwEUUeYPIvZT20L3Rrgy0eAOcvzX0mxAoSgOqUDct
8afVtgfSle6RAsKvgl2FL+QDljdM78WvjfEfH77aslllyK20UcdHgNjQBb79Ba34
9l2E6/kOPQo7J0tRcOHM27beyQ6sRDhkhaBumw5Ubnqgo7C9ycHvJTJU1hv9DybN
CMd/V/Q6IU5Y1rHHCVZewNWaQ917L2LZizfdl2tuHTBRiXqmMyJYGONbWUlZ9AbZ
tj+0gp6t6xsHmRpFnJlIk5C2tZdTqob9zYGIIJjNZe/TOKSk3FsvI9hsUbKF31sE
uEJyti9wjiGnJA38IpAjNtpihRa+UKt4Xr0RCpa8K9ZEnfURisuGMNTLMc5ngMyI
7dfOxSwfNcbtC227NXrvpjT25ZoOOnV3WnToMqcsfL/L/om/eIKoZm7jQALXNeHJ
e3i5okrxKRf8+GASvhl22iSGX87Wwf+oWssw7Kh+5kDpM963/SWk4EFtjaIK5ysD
hpUZspZ7dWaslENAJiB4xgpAB1WtecqYNDwtwUspyggKCZeFFTyFGBUxE7Htctb4
7SfnrNBzCMVXjZxguLzDxWIitTvjAB0FXNH4xO9szm41lH6r9zp3alDt9RVmJrKX
/be7XocN61PQUOQMKTg7yuYyM0+i4GueVshASWnei08ZOq9e0XBF13i7AYZSpSyM
SUuiuaDB4mFBwnd0ioBjK1cLXAcBxdjhMFcPd2Szy5uFOLp8k3XBk9SsxtYWGd7w
Ll54rF1m4lQ9BPTDWLkTdwFX6YJ89WT/zmZoZVsynlOtiE55GqALj4/LpbVO/gaQ
0aue2MgNdP3t5VYbSreKDAu07UBWhCuWGDqr2VTLDeSFbNJAcyVWoRb2/XIingfT
r4cupiUmR0IZTqLWR5y2UDFoAxPg91tJ43IxWD4t1d6Ihp4cjNNjTd4In8Df3GIz
kQf2SJIYB9wFzcX7xUhuYtZsNnF8ZCueq72i61UMoZhOy3n/5VKex/Jaq6XmfMnx
WoVB+ZMDOf4uN4cx0theyxG0c64TCCLDEnNZY889KIzpIc3dBAgF3ylwtfIvq+Ox
YFkgKf+jKuB9Oom2s6WHSal1Mgm08/kc4eQY7rSWucxwzPntw+3jg1EJlG7QlI/R
MXb9wEHlXa9EA9cZuxLZULJx90u303h6n38qaLMD49PJhZl6iB4ZYk3nUQjifuIC
d1RZqXHkLBklSqDgxaqy+XqZSkmecWxal+qDWAlQI8mxVvmJh1zIY59MNLgv/Xf+
UphgzlBfiVHnVXQP/qsMyTnSDkeovXnYAaTHIUWLNJaGAFnhiKA6UW5OJHW5Q3YZ
i5L/n+DRhzo4FahXm5luIMFnFY/OSnIXJb2jFExUfF8SY6i46qUTbncnYg9Llqsg
wNGdAnyNBUTAgBKLg0FY2t7pes/Ylyb7+j7/oz4WNdrYPHcALLE2YXMpxF6vDEkt
Xn64eqhMy2bPFOs7pRPnnWh0eFL5a3WnWzRJbQZAsG44NgANDjkFiKKl2z2emvwU
Xh1P+4E3l/NeOrhuDhEKyO4D7tu4ubKtTJwr9yhzy8XljYqf91WAK5cYdUImHBmT
8kShyKrp8/ByrmbbH7hxxPXv/RbeLsmHmr0nHLrd1KwwzburUjJdz6u1KyhUT4qL
PeIRAycOp6etZUyt/JlTJOolrUJszu49mcb9qzYNR1dai5p4xxn9HOQYNbSULD1/
crKyR+wCmw9+BYGGCr47PmwHTOd1FNF6SB8FB1lO6QAdOVj+3MawcT+HeVkTjHI1
Dup22X7c0dBMfzUEflZjwhElZfg07HxG4bZam8/YU6C7+Jn9MIGMwGmiMoApa8ex
6qFQarGdypdu4YqVP/f426EAsYG4LruMrF0it22jYteAEElag41kT7lDoT3PQH0o
Z5CJT2I5IVp5CoUfSujELZgh9WmsYIkGWpRC32NFaYBGsrL/vY6wZUsFZ7+48zrg
qESHtfjhpchzjaXFz0prBYG3OvoGEkCGnOsMItq4K3q6PKyLG3klU3ENOt2I2SSe
NY+rE+P/Gr7NXg+9/zCLJiaoKAO5/pnr2pf79dPzvzFv+bFRKga/qd9p4fZQ7HVf
iUXzylfOap2zmCLvTqYgmSlmSjudOR5902LbcwX0MuXMwE5wdqchWWXquFM0JYLA
72dDaehT4TJUFNf3sFlPst0ItSuYC01UJHPhtNezkkr3BiN0aU2Y+2FB2ALQpM9p
B0/1gN5sZDbf7dWwZIqSoZhgYiY99SQPN9e8+HG7t5LGAL4wc1V7EpTfgwVx0RCt
tkBY1Df9Pf8r0MsQgebiekI9CQNVXOPCwDkU4eKtJ9zcHykw/ARt6eMsw9fTU5B3
/YW7AnG7sHzfl7Whtz+rkBCZpL61wvGQ2eXpFMi+U1KKx8LdPSkov/+4TlHi22m3
peO1l+gUfVZLz1AsmyRhpJTB8TsXhgXUVJf/uTvnWFvT5eU3TbWmzQ7y6SCpjTvp
ac5RB06bVwpM04UYhAImOhrEfAF2m01+vqZz7s1fTuBTdDEiYqeHlOt9woYow+RY
RxtwJPgq1A4HIes2Dqc/4Gq0RC5iXj1Cm4ls/vi4z4/9koizRv1o3zv4vy56J91k
NG5d0SmPFcMUAexP7DzVIDibcu3I6hI0isPWaxG0DLKFHNBitEyl8i9hwvBZX6SL
1flbo8I24NB5euzIJ6BS6UxobFlYuiCjs3FLP/+hZ2kskyxdimo7yqnNNyvraaIJ
WqxHe8EebMwGnyHO/vjtzwZpEgAHuX2rFJLhtycoxFxG97N68sd+Y6rUeGtukCWz
aVY+VdnhNO+rQL2UaFsN1Vme6ow+21VSQYsQKdseMis69Y9pZJ/eqindv1wGnLZ7
CpZ6RtQYF8t4i8+gKLdcp6Tm+/hxjxeCxmSPxDb/em8qCPDj4k7dmlgrmRMTUpcj
FD0KDN/CR7jamKAECZWYj/HfX4IBWuCgGxSk6iMt8EJ/GCjWvMMpeMazog+rOCZE
bJQNeEs+teb+OoaeyNbGmt6LcE09xSLMKfk2d4/GxqbHB0UViziIx34Bacx0/6vy
QqJ7jqrpfN7F7zIsqQ/KZF/3SmAbZRxwUzf6MBaOsG+dueXVabwDfYrPK5qZh7Uk
ZyvMcdrm+ACokLaa0PK2QvJh3BLU5/SXxY9dLUoArTheuQnAhduxdCCzyuY493VI
+1DmpKY58zNEtKoYwrXuUwgoaXtvCWDoqi+W+7rtBOOOUBaszBF6ggUh6qI7AUNS
XZ9m1UD4cH+d6v6r/GKgiIrGMK+9h6L5jST7L6/BhSoW9gS2DaTsWLTu4u0sqE+Q
onsRBt7PxPZmWi7/jjaUT0NoF1wZRzRwcRrHlxm9mSkmz4qSIrE6M1zBrOeh06jC
lxFtUm8tPsCoVGRoEBj8NOiGHZ2zNJOIpOUCwj91UwkA/SoPUWFbcbNikm/6NY5l
oDbizYDOV6v20u4eaYkzxnrLUEAheQQllXemCKpgLSYqbnMEV732ddFgPOC369g8
qO5C23b7KFPGIcd/5OUAw3Azp3ouMj/P5CA6typKVFe4DX4q9Oxf7ihz57JgAnQl
vw+3HlH20TOqolQXn1Fe4HQe9YKwCOCgN3Q03eKcBroPeIw4W00Xbw30yVd6BwZ7
9Okef+fTn1AvD/uMJ/6NDI10xoOjhSUfq2g0x0JFpVHt76sn+dPdj59GMKuhV4y+
MXA6tvB5RmK52N4v87y43baFmZCWJVPA0Rhv0dN9erWHtqxpVXltu0ImvYDywoM4
FkYubGo7gsE8X0Snk6Q9wCq4dcclNAlrDpaRjGTBoiO2RzjphNr9e8aItCF9F/ud
Ui5f8RTHdVnX4pO3Rx27SzL0v65Olagjahr8OjyPOJU3kfqgIWsCUBIwdoMralcr
CsNz4IiDPWmO6L49iFV4TXTc03W0ttCz+RloW7lSA840BVtPidRxI8VzurH2OE6e
6Yx5/qtLuM14DBG+IKKghKIMqwsbBJOmW0dedxmDLwdNS/KNKN3E3hmI66176hIp
PO4ZX12Ka8ZtEQxyNY9y3C11rSJAYwhJpB/M4FgikH/LbRZ/YF0Bl9meI9U9hEWk
RF0yr54MhRNFfGXY/e9F9rED380qH4Gn9gTi73NUZ5MIi3wP9yRS7X77lFk4EDtU
rbqksQWFYV+K6Ia83Jtisy99495UyXNWcfihdZQBTvQdm5iLwiGBDAw9RHU4aK92
0Xl3tlhQ7MpnWwU3SV2YlYoQcu34RCAFlhRcAfK45fJpDuiSbDvOiDLJObUhfd9e
jBO5Jp8aSAtCbhzoHOrlKq+adzqowgYhh5gPoH0cFQscFJWwc77++JIjDzYR1jMu
OBN3NskoxutJtKyt7tGP4GIfhSdccgK3CnKJGxlMcasrKPxcZ6+cvbrgwaxjZewU
azxyS8X/sAGA2nd0YkZBEmV7zHD95DRyMH+UovDeTBr1B6qYUXaxZcsMNDxvRv3z
WWf+kQz8NAcX5YYb3iOan0MZtiQ/6vJhZ9HBz2+3rOntcPUsOB7zaX+7PXGAskhn
dQ1lkoTwEHAJHHMPCW92wyZ7FWnKxCUWThZmun4e3ow4bNd1AGSUOJy9sUbx6gKC
j2ivi74F1qrIpubuEw0eQszfEJAHc9S+X1T4T+Mny57M1V0QTg7RmUJXum97owhN
8ykQd72Kq7CPVrIwGnC4Pd6HbRSfcL03wYRFiBpE4+UZBLgcPXyZlWtRm4jvLk/B
QOv1E3gdE+SpBG5VNcWVFBFS7aUDoolvP9vaI/dDxX6yHPmZ3vCiOnUQU8MgDMLT
G2ULfvUL/YJNcgTwU9uLlriltVsebh2wV0dIU8VfCAekQRs9rLWzCaEIhkN8TTeq
mGGqIe3EYhRR26OLFOTbyvpBqXSGz9eaoogaszrG5ZoaGDCbYSUBBOxkUFbxWx/O
QX2gg5QVWmE2Z6OIcbUu2JiHaG7QdCyVgX8NU9LgbjAuRMbfMKGaTyM9oXab8NmP
qUeNhYyw8PagoBSrdVqQnRNrv3B56C6Mr9mGA70okeR2xA9d78oRMv3gKt85kJdn
PVOKXp13m3+j45hV//1nDHYiroY1bY+Hj64wfp1d026ayMEIqU3ZG2jSQtHxgS6S
S2ApNWGJvFtvEVKHW5cRUZWSsgNtel1CNuZyySpi5z/BHoHqUZ50VqWlRkI7lZxG
nxvt37hUofDdaIvmHZgpB04gjYND9CVQrSlT5dYmWmV4O+8eSSLwxRCBaeoGCTs4
kwey7iRLS9R0qhOWJxi7vojUj+GnGgIgelG6R11Su3SSjAlaod0sYESkV/9DKbl9
1VJ0O/pVAKcCa9aXZhDYA8lL5EKWfXA8zWaqn7ls5M3zxTJWto216i60LBR2yQ4N
G/IEHD/5VDsZiebg970jCkAMklEL8CaxWSmJeIsgijgtKE9tFMwWm4/hGk6U1Fc5
k7RvhX8lj5ddQat66c0OmYynwCMiKrh22RywNEW8ATGtulQF39+y81HgCIa9D+Rc
fUJvIKcDY0He3LXEZU7q1nMDNTgam2PWf2TQTm3oDLvT2k8+xn0HBGz2sHWrTKUo
+eS11D+ZNCMUcF6iJp4Wycong9KyqlnHYa9y3+shs13vb9yZrNcUszgC8Uo2TWxc
jB9qU+wi0U8c10nrDQ63k4aiRT+PFr27A09JC97AL6N3AkRmBT1I5awiEz2pKc+V
VMeeKs4D17P2+GSKdEODK9Wt3DmpXnoys83HwZmiO0+8ZA9vMLdtc60RXDDQi1CA
26EPAvZhw2thwVRhaL5aAMGmO2aweUwtvzwuaJKno8sEUpxxzZyycp1qqsJ5aV3q
0IPm8nsNXDubOZwYBtAhxCRzSdEE6ATJa68ripObt/E0q3E+0A6XMh+QxW80JaOW
uXwEdj+0WWHwhrquPldcFMyv2EemABQq/Jnpg92ljBOjhR3CIA5jf46qvYwttwRM
u4vcDKKV5rDEp0CWBM7w03YioM+6yZKAVIspB/HVPuJxX6tqKpvJ1pgBthGJkLvs
1H+JT8VrAdYAsaKCVNIImJVOSGnfL7zuA41pfQY+GhQqxsCpf+OhQWnvrphEHCIQ
YWPxfLli82CBgSwhakjTW4Qgvy0zPHfeAmErnyOr9WzO56ZhCT6ca47Nx5eZL+oy
dW+yRBb0z8QUNbKSqASX4e90VKymwNX42ldgNh/1+aZsbLX1gVcLfuTJnPgNdGp4
n13HsoBczIrpV+PUXRsEE6ZnVhLn9abckxt3MSK7DR0CNksavTldDda/5wF2MbWz
P1x8qZ7u974Il9rftXFyDqVSlM5aAlp/JxruzUUCw+6xsxeFtzlwZmnLCcMzWmRs
FiWZcuQ2nVZv/383POx5J2ochEp9rVPM3S3R1gx5R2C3Q4GfDAnf4AvZWZW097fp
kW8S6x/Ht7JGYylkEcfe6mrnxr/w+Sxzs2+bk8529riI237Fd9D5fVNjxO7x6LLC
K+9Y/QxbDzv6iYMNZ5DsgaxT35TgWdQIEPYzxcqexJgq7bGY8J7+fRv9GtCijLw2
wNPLU1zgzOxU7x4sYOI1jwEgW8mXoE0+cZFyxEjdmLkNAbFl1RPYCXRiuCtZY8gw
oZd/dEgTIJefY1/GpQmBfDLsqilSWaCHFZlD+v4Zn37Af0mQZeDUDPmMzocpo9vr
WUERncbKbG5ZHGQHlIHtrB35K9ApZGpVEPmDEzNGA/CmPOTPPWIS0PBUm+RecX1u
sl92xzZhJMDruCKnuh/EUeQCVf4FpNiRv2HJ6h1XZNBVbKhOw5J63S+oYn3DLD2T
i/RKTUu3rIKrzj6tDvJaISOwseMD1sbGDUSaUZm/BNSEIJv59+dKrKT42pO0hR6E
VsKc5dwT4L2ZioPKvqBntWwc25OztN9XqDhHcn1ei48cRbPPhCI0EhquSjCHUe71
5I1ZGtV288ixTc83CxN3emz9kZ5ZQ6/5h0WjwJrqUpeY41KwuhL+Sglu1/EgQYO5
cHXynuOVfLr1Z7U8bJPj4GPxm2XGJEwG19lPNXTz4PWUPp35OvWg2cy3+lhLdPv8
94pJvZoAi+U/Pg07dBH71ba8rMQbadqqmJMw8741j5ACLRfSvaycgQT/orbBBeHW
6zI7i0sfOM2oYuGOpT8FXX6opwax5lswrF4WXQVtPzQ=
`protect end_protected
