-------------------------------------------------------------------------------
-- HEIG-VD, Haute Ecole d'Ingenierie et de Gestion du canton de Vaud
-- Institut REDS, Reconfigurable & Embedded Digital Systems
--
-- Fichier      : avalon_computer.vhd
--
-- Description  : Sequential calculator on an avalon MM slave
--
-- Auteur       : L. Fournier
-- Date         : 19.08.2022
-- Version      : 1.0
--
-- Utilisé dans : Laboratoire de VSE
--
--| Modifications |------------------------------------------------------------
-- Version   Auteur      Date               Description
-- 1.0       LFR         see header         First version.
-- 1.1       LFR         13.10.2022         Correct behavior readdatavalid
-------------------------------------------------------------------------------

--| Library |------------------------------------------------------------------
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
-------------------------------------------------------------------------------

--| Entity |-------------------------------------------------------------------
entity avalon_computer is
    generic (
        N        : integer range 0 to 32 := 3;
        ADDRSIZE : integer range 3 to 16 := 3;
        DATASIZE : integer range 1 to 16 := 16;
        ERRNO    : integer range 0 to 10  := 0
    );
    port (
        clk_i           : in  std_logic;
        rst_i           : in  std_logic;
        address_i       : in  std_logic_vector(ADDRSIZE-1 downto 0);
        byteenable_i    : in  std_logic_vector(1 downto 0);
        read_i          : in  std_logic;
        write_i         : in  std_logic;
        waitrequest_o   : out std_logic;
        readdatavalid_o : out std_logic;
        readdata_o      : out std_logic_vector(15 downto 0);
        writedata_i     : in  std_logic_vector(15 downto 0)
    );
end avalon_computer;
-------------------------------------------------------------------------------

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1_1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
kD9mq6NJ77uwdpvfr+ivMussMxEqJB2Voh+X6SmuwbXYEbhKwY8ROM3+3BCoEZYX
sRjqbKesqFbFvlOYjqoSzE7yVsoerOH06qEEpQCzrTu9ofhxunezb3jJ03aHtIAV
YX9zuO7l6D42zEPfrK7W/LbpGKUGIPjDIe2AZQTpleDVxjQHLbkRPb1d4SOi+6Ej
RDWXCbAxQQMnb1jKSPWk+zhBTh7+F4JVxZlbfWLN88dD4JJCfPmUtaGfbDD2DfWJ
0M+EB1AIDxmKb1/E4jUGWcvcJ/lBKknbID78HVLMEGNODwMhamHCoNOx2dG3uz+I
9rG87baAj4LDWfC9GVpr5A==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 20432 )
`protect data_block
r9cK/YGwhjMdBijO5JU2g2ZPKcxJN99ByA5t3hdXC+YMFSXQkEsDj8TE/B2Ky3X8
+wWNDlErLMF0F6enpCq9viAdIgraxEcN4bn9cnd7yehGGD+p3w0cKfUiCZ62KoFZ
C0pInR8OzX/cWuHY1xsaLRLjFtjbi3Q9ZIFPBIIpI+uZq9+cQ5V/BSWZO0L5Rmwi
kmAXTRfnrLy4xqPTe2X11G74w34sGWDfyh6u/2wzOsDAeUtQhKnHArGWy1JfAXEb
LMaFgvIID7lowwD3d8uJHEawcymJwKPNgGA5FkJAtBVyhBeIvb5mvBorYoH76RoJ
489L9O8tmEDBnWmwbIXSol6OONwJfhQwPHi4M0zeE1ZNOncDWvvLMvnz2Yox144l
QMfbF/zosZ4Eqmp63aqGFplxRnxnhZAyBnIy+UBNyICXL5WPhbW6kHVyS2dEROuP
id17A8lE/sgVkxcs1iflGgmHV4I1M7irH7tgGjjY3itYwdPIYCJlXxx8avvMtDPX
+L5wax7HrOg3mMbluLy35S/FmG1hwu92925H4OZq8s1NP/E13FQUzhLwPYBxeTNJ
ZXA07YwpP5vBqrOFpoqjQymFZ2VJPvQYOzYlhLzXIlqg18a75ldSr7+dTYMrd79m
I78w0p/I4/IO/zElI8HVurnhLQVn0YoIGwYOeL2f3NEwJj/SEF5XSOy9mXxnZ8rP
pd1y/uakMzvZ6bqLOl3a29ga2k8OyVljXr/p++iZXQz3XDkb9EWVpKCtjSwUvOoK
8P1Bh/KFUeth3BzVotriP0EjnxDEP6Llr/vQsRcypR6fjsPN1KKTSWomIzPG86O/
0l5m/1wsoGs4oAbNak+Hj+lS9GDu53utDVxX7DaJvClvkDwGGfJVTIxyHtrD5ANK
HyxRLE+LB+YWSUxNVU9aRotVbjar/Pp3rsUPcDpZB2dC5N5dPQih4OZ9P8HFgK1n
wkgRSM2TyP/HQ2bZEbs/zblbKwlWzOwvDSwcdD9QJZtqwnD+ThJNi4nVLUTOsPw/
esdzJkQUI6g8SvAJj0eoPwXrADswQcbwv/WqZyZyI0+W0lTdXqB4L0ZOO7+XYR6w
EaBMQkX5GXgfp/s6rkqj3rCjFqV6EvLxD6H8D8yvSgZK1MvQG7i8X/1mZGn7C9Cv
RAYyiTuzKksXRejm703tJTRPWUHxIJZYfe5Avc9e2nDI0VQck/uJOwZPH4M5zu8g
CYj5u6GCG63FPsLBUkGgaskUUQWXTgY5Jbw+pB5AvAs4gqDZZoOB/hflINbY+keu
l2sT8gKVKJyNjeCntMJGGglKL+h+tywatu16XcCgQgOhAJlpHjNb554OnLhatV71
WnFhlVDyxzi9e+DPBE929rqaAaX6/B1PTCz1iT9QokoG2myRb6qe4MA9gGBNA2mx
k3vMh0rNtl5B7XXbPMMz67NuoLmgItBHvDu/X6nKhQgTLDm74LLsC5BCVXP6l+Mf
BYENjgfK5qhU4ur8GK2jvwCNh104k46VF/Cs6yVO3KGBQQl7pm8xvZOsTVUSvB+i
706JuYMDxvDvhKslB7tkv33S/RQPcpiHXRpxrSRs9JpZ/ASQdwl9N5nxB8t9WIm7
Ssbbxl6XrQvMn/rphMd/FwC+GcEZJL9yWEbuj/CgAmu+ZMjFyuvyWA94BHgA29mb
tmSESHDrGBBc8nV60NXtRXlGHWJYtXYxQaZBt6a4chAlF4x9IaVn9nASNMGZL5HX
W+TBky2RyAQ43IDmrjmsC8u6SniVdSZ+fGTfMTSxf1ncvdB/xrwtJx+Ozx573RAU
T/bQTTAjSSejyGQrp6TcUoVrgv8uoJAWy2EC1Ece/u1lMmQ9HuXfDlGKtPZITJnP
0wjsLpW+atm5xaTct8Spbql88rrOlZUfsil6L8H5/EdAhluGZ6sa2HsmwnFtmw1f
oPeYBKV5OOx259f1XmV6UdyDeCM8khvOFYIihoXyVWFk4dCwfDB5l9PBSWgXeIqk
Wo3T7Q0ohjiMnGyITb8BV5DfqTw2Odef4B08HL6qq94UJRjSxZ/gPI45O7oZC8NE
lgUu+CAF/STpnrSmIddBAjK9qO+LGuwcrOXT8WWs4/rP2UyJZyqsfTDeNEsENi0y
Sswf0lYeB95qyZChyO4ZO4V3SGLc8RR/ntlk9nPYbz5eHf+DhWWLobAmMP9hQMJJ
i52DjojAc0euwTAcJPeiNs/pTaUcAZotTIS0ELLXjKu7bsxSAGLsjUrlRjX+d1sU
/Hfoon/2A0aXOTtmWomuCm+/4Sg/E4bq4xe3nxK5DtEaTMiN4/1deEsQ8Rjg+MLW
bF/2SJixJCcTNQvIpjnp3fz7uhe3z4lVBwp9I+GMju0v9G3LlH1+EJ09GJA5KY4T
1kkTSsxYaGefS3zn866cBwRtihF/6+F5gJwZ0xHiWyi3M67f7gdpPzuQxJUndUer
4MlusyAuTv5ENZrvdw0Cz0Et0CPSDa67omVvyeoL8PKCXRgi2U+ppEFGr/aoLnIu
s5uQ0oA9xi9fGyc5klCxVb/o6FM60P3CHicaiuQDAP86zKM8DpyFMV35RooNWBNs
4KpFnRbrn8R9ytIEL+P/+BaE0tUq0g/6lBx33TEj1lTTiWkU0IDXligzNk82n8pW
vCWMmQd1XQlKThb9+8HKq3fPRT16jmOmlt81nPTB3BudR6eKa9NcKwcR+sKXz8Z7
9kVnihlWLpVpw+j/wtOVHGy4uzb9wB+/BV7kkdGN3tkqF7z5Tk7E1HbhjsctjkSq
R3OmHG4wrzf53Fqc4XKOxvtcMFbF4Zkg+PDchgji+2BXNAj0M5LAlRl1xZbbTI8K
9hSuafcEpETzD3fPjLgpyTshlbj2z82PUdNC1gEfBbYnzmXOs2s3xFdTgTJ1mKyR
9o3MWb2h3dNEsA8EH4NdidXeW9GTJw8uJaVSu49RTfE3ceyRzZdVWWP2ZVzf4RCH
iSlCTOjPtycUF4Kb68Jm5+3jc++x0WffSbfE52mmhDIHXkEYhlcCPwPwNS3nEv2Y
3pl42Tj2SB6rk1wT9JZBpEcW/XkFFMuawEW3A+MPIKJLYj+QqA+icf0Lei/4Yd37
zk4wWozMEFJMsXe8fT+diM9GIhisMve6KI1QQuw0fAVlsy6ymi/GJOAY4HSVJuGo
jGkOBZVKthO7q15ICdk/W2Obzp3O6Gab2Q7+FjtCm2fRivfg22u82KBJioYfv8X3
LLuL21FTvecvozX2lkD/ibk39FAgzu16kzioFhukXPfxKv99IaowE0gfsJrQYkcv
dqQOecB7XooLd6DrQdSwUQtqaRIfeR8zFoeUNdrELX+D2fUDuF5gu4H5/AVZe9y8
68VTqRsInwzZsXWHvKi3+IHKPcFEbWj24RryuBjuUxAfrPmqIZFQ5NETNLvuocsZ
557Iv9HFR8obrMcT5W21Fa6Gor1I+mdkoHJ42tGaCDtaSm1py7RGhvOpHGpAJxOE
WXA3oYVvruPWMZ+hzdqEOKfRFF72J35gw9IkWyq0XoIrNgHCOym80UNoRvLcYaSB
Bqpy/XN1mHR24N/YStEziQpDT/+xO7jgNkrUIR//gdTGranIgHS8gQCYLX18owp7
K/4DVEYT1E2r1zdcQxSqwhN+0Xat6nfRA88i10b1n/uVvv0dTbNjPd+otcLi1SeC
dp0PeYBgKySzEygZR2X3MhgzXl4C2efyZAUQFReCw4PWS/7ybbceVHRt2HEdBRiV
4Jx3Ei7p8Gr2UbCulUQvB+9fjyPHnWcXy3tPp9Gbrycu06JUJfHGTxavIaXGyzyO
7s0J1x3S1J0NTV3bLbYdPvswxJJYawm+JwYQylOAq50BBZzfJbeqQilVALJJ5LyC
yC2GWMnp9FoZ5F/zkie7zCwvYC630i6xAVYrb9Q8SZJ73+4iyxMQBeMi4G+Nvk+Y
3Bb9PWyKNO4zHb4mvErNuuknvLdOOLYssazC6Pbn5+zGCGOndJBmw2bh1bp6/0zl
pMOtmFs++vQhr3PDdDZ8P3ipIrOSJqF7G2X7o2p+5IN7IB7tEqPLBd7F6iU7zxbT
fpY8hcJEYYguZhrxRO8cUt5wUJGpbgatJfjN3+CCV/2wlssb+rRn9T6I7bP10QLg
TI7vGEqTW4WKrMyOQWifEDQujCp3magYjvHsQ6gpJEC0GL8on4qx5Y1PoJqOw+IE
xnNiu2PKrplyY0MxZwsP1eoz2wTBN3fLGxqjqucNxPSXoI3yt7KqUQ7n88HG2GwL
8+0goJlbtbIhqRQODXyZ0pXS0MpJUBdH7qgbo+d4lr0V6/j51tYmLRNkjOcmD9i8
W83JvB7byvGn9v4NVIPhFcg/iXztBB7XqYLivxnJXGmdr4SCd8hvm6CU8Jw07VtZ
K6aivDzvIgptVLKL0W1nHpoeK159CXGfGxhCosd3rRNDXqFkdv4untGfFqgQG7K6
lT6jPE8eSysUpdVeVP24khYFfyHqske2/RQp3eA/yYhKkad4IIbFXJwhK9XjLzUa
gVNR9VKyYMnZff1Hf9LqtsS1jiZJWEo6v4Qps/YkHWN42jrvBHHZ7tHGbNlavLKu
T40efEZGKhCtBPsbKLFqiAX9sDEML7UI0/25uJgVxEwu/NlryiwHS0YQRO+yz8fI
kBYPeanS1qrg9cnArx3B7eRe5c9cTl/UZ1NeMSz/LLIOBENDR41moynOQX2cyPsr
mDbrj6s1uLwKROdVP15K38FEGtvrz/4tasBwoRu0C4w6qmBuu3Cl9VnR8J9ervk7
HYvbdgA67HNna/bgPI2NtqjFxbRWKpDXcEtgDCertzUli+a4iW4cW1rI5ymE7pMr
vyr7PuZMtWlPuXlhqe9rO4IkdoQv1FbNo2ecahClQCdmKZaOYVSaTP86z2cB/WoE
KOzabr9iN7VweW5PaHm3cCmi4MPmOSc6HCU6iDWkRAKr5uP+6mHqVPAwjbwIx4a/
hM8ENJdsX1Gwl6cgC4b6ILtaqvCedguRRekumMBvVa8bc3pe5pORGf8nCljhRuzb
pc2N8BWgwEBehIVqq5zuA5aECmCxzwKVzlB+qU9UAIyMnbMDC68u2vvRkpQ3PogO
W/lyaA/WleZoUHZCjVPjzp9qHXR8wYPgR5KOKADGOVb57kp/i+maxhxqiP8kl+h7
jlMM2YxvY4WG7Jqp1RIMIvwb+bsiqO9MTIegbwqULvCJl2AHLXS7F016fG93HQnx
LVCTgYKb10ya+cd5ifCAuO/I7ko2AwaySSE1dPqC9qqBnrMQoe5NhYdEdIciEjAc
A+KID+xugfCC1vI6M8Le+v8Rw1av7GQa+aWgc6D8kaB886rAXFEyqvxTA7xOsELB
21IlpZa7J07LKxNiONqO9nUkkAQ+Q765yx2DCwjR1Y47mAhmZlIhA/PM8pGNYZ+e
vpHId6wjdlvxsSEtP/WAVl6klBPM/G99xzgx7kUuOCCICTmrliPIJcln9rie4Nw1
c3wDPLm/45nnt2xea1cudicJ9gihYQpD+DCF0xpvX0sTvs/TSWn0fgT5RgxNgUYl
1nZxUUXI2QPiJa9hG8p0D+6WUkM6nyPuY+AkYP+DKV3I3bRP0t+tBHzJwhGxxthC
UwxW2yC8lUQjEJJCVWPrBcKeLIio9hHMYS9DS1iqXqdr2SXiqPaH9wqK5CM2Blu2
D3wSyC4i2kHapjQucyT4ZsNaAsUXTS4O9g9ksI3M8nbiooZ/JBAexiuEik1sCqvT
Qh6P3uC28Y67u1TZLc1CzscjVxO2MxT6frCDWdzsY2+yPrMd/LVVvitCGlJTRORY
26pcAxRu9zVUxmjIC7wS+QJhmGdPrynyMiO+OmcBe5rTmfN7bJiyTW1Cz1wjmiH1
9chezWyHq5TxxG5R12zlafvosHyyFP24H2pAGddexIA/5HEcydFJfVCXHV2xZBLq
hcBVQb1i0Wy/iG+8Acwy+A0uxsGaf4YIn/woTgijGs2aVZHrhFZGsQa10do9zQlG
5ERfqkRaJdcXDywLt7fWd37AERpCR7EWkyNy17+PzpLGxMFYgl0vbEpHUUJ6yXVP
1u9GTMX1hFCzsZFqa9sOsY6huo3ZXDpZoibDeLryrGo6deH1S9V5dwtGIe125XLN
zI/3hhOStF3N8VgCIPYghfYnVTc0sEmB/7iHTyLPLBMWC0nyFJePb/iYtszUnpwK
RbXJh30uXuQLwrhqk5UM819iWleIJYnFmj5XXKzzV1MFcZZN7WCKlPYSR8b08PkA
NudzzF/u0MahE9oaVqG0HqJ3om7aPyIMckonSGGll6lDxAOR6akgXjeJ20yK+eZz
cazGgzS2ioQw9DOxe6k9Qm0RvcLgZFG/6Mg40R5ILjJErGTvSwvZAq8up5Y+I2Mp
BQaJlKrLFTnVtdWFQKnUDrVVtbq/pMfPWFIJDRSL2gIuQxSf0JJ730k1LuFA9bK+
N9bTNSi1T9jVJjm9J1F5yJxUtsIQwXopu1TYLc61Q4I+PDDl+nTs9eqUTr620IfF
EjI5kooPyYrw4Xuzhe2HnTEM6nyP9fuClfIQLlfu+LfqomPGgVyTIsD0wJdqjwTu
e7pz01VZIHtMnXYPRjJJ1LVa5lfkBpMdxItYX+DLJTpLEnSscfiTccTsifkAoq1F
/lqK4JCX1naPNHRwAPq2qiDAcHYSW77XOxOyCucQCoNVQhx7cGNpGFoeLC0HhX3F
+bpZQAU+c0hlIwqwYybEka2291gcimVJxs3i1d+plDIJWInEUeAxq8B6gNiXX9Fg
fvg8gk7PTWNl9xtykjfJIYOZGuvq1hXctnfLXlMB2AuGGMPV8TN/8NB+xpfWJlym
oN/WXosjb/Jzws7eYQOpDGNZKuwG0Ak+LtMSb++PKPkECLMUY3UifVFwLzOhODOT
hIUJSiDrWxKi5U7ecDVklcKFaotBmiz+J2Tj6v9Y3la0UwXvR/A9V/jJinU/rvO6
EYMUcWNDRskzCB1B5+IpYim5ZC6RJHLZg06DeW++wLzCbJeAzR+iurycNrZIrGkf
TYzKJe1Vu+7FFaDMPFLebP7ErrdQQSKCiS1UD7OuBilgnrZ5GS5lj+HHBjTk2pvx
/JQ81DBrEHRyTD7YCxlxqr9gWcHyD26gX5SGHhHzBglsS5lrfbpQn2Fx5UAbREG7
uVui67s/XwCHKTjiltQBmkg+3gtHjCeVbLYw6vcuBCxagURXdxgm68BhnBmo37Ox
PcVFq5/6LyKzSOEuXJsp4CXAij7jxVMx7g+2CUrvEqc85JwWUEQjJ8qdpRevurWN
gjIzlXCm+t2ExTlshs2dkPoAEsUyN/8sr66A2CxPIWWnzA3BfwtFqWI408LLVWKq
Qmc08i15P6lVyXve9F0UGwIzOexEXMMCpvTI/TJ/9xTCBNwsM/QbkXlh+INjh695
c5FbqUF57egh+TM7BFO0ALfbcDHdNGXQZ6wGT04VZSVK1fBJJtKXcA60DUPY4Kxc
LshR1xfHsy7UPx0DNLDhDmkluc5K2a6cRPDHHLghp7ORrVn7LRl5Aq7xIMlHytuK
8747k8boYS1/e1axYmhZW0RcwVPSjbeSrj81TBNzcAUFkP99Aui/ZmfyPOxP4ckI
8lPiXq1q9mBGsCxJALn575nzcBA+JmVyKRdG1RrEAKXnu3mdRW7L+vP2g3tHo2YP
x2aOqJD27bVrmMxz3UtMNzrm7dDIsOfDRWiR4leFJAaWUgRY0lRhjWZsEScwxHl5
t6ulsGhALgwW99ag6Rhnwmc3RzFsjqIUeHnfyDqp1T72h/hwpACoQ/bAtGs6aruI
5xhBgfQZIBqMwFgJSfIpX4bpVhj69Aataf2ie2znMpCg7NS5T3Me86PbreplnRvj
O8HAI5MPzZ6cTioP756jtnHJIlxUAVyxOrpathmR5o4s2mijB9w6QAR9Lxxef4ti
8y32JNXI+nLuRSJwW5Sm18TEG4Vtr/vG4BDanL1PH6Vsofwt1QgWUYa/zAE6L2rM
wfw2iETsmuQFTiIMano5r7HViaEtUEKCyzpyeqBk7oBKYRtaKPjutUP1Br932cen
IZwuATMfYT1vDGBA+GqqwV7Zgo5VsyQ/2F++R6Vb39nwPq2IFkxkfbeNkpIJI7Ip
8BCoh3qsb3zoGwSIo9Nsnd4YiAWpUqKy1U200z+Ov088j4iBHtNUu3C3kWnRO2/U
4x4nloYTWkZ+WJZusirsqbagtTxVWTgHNO8UgUBYMTpYbJgr9AOOR7OBke7S0gs0
PddKfSncrMm7f70oNW42FSA7/hTlh7m77Bh1gIoEPrMTOj5WMMseeO45lMCZNddK
+2+YLf4yGvq9E+bEozU4uJhT8G+yJTF09GLdPau3yezhxRRzERABcmWtLzSK7rWQ
wcN46VbLKUH0rt/avj6FU00LWNLWnGP6SyRvlCs1lC2nNoVr2DOYVIsaGBhSfqkC
EjFB0PEzQbBpwdB1yMx9rVQ5CflzzhBqkpPP7Wuaw290r9Uv/6vKEmtrhvGmkRWS
yiHqCmlNPNLy1b63syUxV+T6I/J4WpnS4+/sPUQ2e6jBry4C9R7HyT1f7bMJUWF1
UWmE7GUM9i/TYblShzirK2t1w00m0vz4xSA61KdQq+y+V7iCIh3gDsLbzszJFL/y
28ZOVkAj0zDDBjh8dHyx6bRog+mtP8UQFCqSoMsRHxpYz/im88hKXvucSfz3c4U4
dLwVYQ+P3GVNo8h9fGRcoBMnpLwv8QGIwv6Rt2Xe59LPWqzoTtnKAE7dh++tF876
ZEmZASvJcfSPNRHgwIFnsl5HWQ/+yAtIUqb9bJ7ZJnh6yG9lq1mkKxDGsr2ouNAE
chCcm7sMOHCihG1WAsCRXCLdHa2DsDwehA+ja3B8D7lnl9J/jwjz5Qi04Gg/Z6xL
xjO8l3bT3Hp8CgY5W/Ubd9J6CWphUaWr/9T6KqH0mcRAtK18JLqWMkjF3nogAF7A
nVj+kEnE7ggVXEoEHrpNFBTah5XTWSmKm/1S0WJ9pN45DrFwagw9nRN68V/58HLe
CRZFXgTZvUlvkPrnI6lgkp3Re7tBMJhctG59WIAQCGFaepPr5NA87Wb31PYkeHBB
TgU3oJEZtU7Q6LDY64moIg5GwkYqS5K2M6PRnssHFLaqn8UP+3dIpGRZbWH0Htbe
yeK/NvalyJspKwBC5r9sb202RQMfeHEw3dTN2ashpm6uFGQ4yH072nvlzf13GYQK
DvvUYgBZNvj6D7eA8m16NSXR9d+wExW3fUzHb1ctz5xwCtVIsAoAq7Ug0TAtOAcx
vvmzT2RYAvI46H1dpn/w3Rxh1s5QuJ/kE9OAPXRercLH9L5ByVmX7QP6z9YyE7HP
5vojq/h4hje16YPTEmAM7qeRdwoseDMEHCxsAQTdrlZcOovcg7Tx0q01I4cNGzHs
EDZOYfWlpc1hFrLp7k9ltcEpBRx/7TYGDDsKSGpzRG0Czvp5hHupUFaGu/O6+If1
kSNAnR/O4VRFIo1BO7YoFq4lEGvUk2WbyEMXDO7gwkJQUhah25PRd47Fad2gTG2p
AA4oS9MI2NizG5eho0iKoWc86fTH1uni+7Ox4sfqGKLYq3whShemDoyD3IJNjGOz
+EYzz2MS+5hH+0Iku7w47SbNe6mccABbwjqmp6MS5P36Ifcy33IuK906a87oR36N
eVoaLD9U1jUrkP5rVHC/PNNHuqm6ToOAyM+DOCOqb6gIYhr0nFgADfBsW3mUnJLL
+6AxMD4/y826runjF0+SNiROSLNsiW073d8KjHX/EuYVxFFjlIqrW3jUOt5astvo
PUUsuX3WAJTBqU0za11sI3xceytiIoku7LXgw+Z7huvHm0ONvz0MbBdVdCnN4W5c
2hjNbR65XpCcTIuuNVE3MWshwsg89WMlYq3Qgv+bKZicrbc+ocX39zjWEwh6xcDi
YpXO7UxMobYALRlNBwmVO0gYO4C7Jz/rWr8gOjzFI8RfhWaYuMI3oLX12PvtWCuS
VjZUcGoOxlvbmhL9Q1Z3IZFrFBoFEKs6O+h2gHTlyW7UH6L8I2XpGIwFGJ1K4NZt
7mnaLqzLCcILuhpIVPC2myty/wjTFQPXKEl4DzMoQjM0jGbtdsWDgZ9OZACBqrwY
83HdBMUNeGGjtOo8TfDgJ6wrkofjI9tU+D7gJdnlmWiAw5gJQMYR6s0Cy3WPkUS2
h4b2Mdy2QxXjwEAYkIHN/uCr7XDuyyQ6Xn2zP2Wi/6SOaZ+I0qt5+KcKdeTpIy1N
p92Qt9gYPUK1t91NrgyKVcvA1VrI1HzdYEtFRjnn0GKFdVhHz3fZbVuqtEvAPbIL
pvkhepCeFB9GZZHKcwExe/ePfBRlcQmwQg4TFcdT++Msv3v9ecbiBRZsVOY0UXNn
q4lZGUsnXSF0GxglBcsPejpMwdSP4mXquQidQOYzuM1sTAIiFTrkH1f7Y3m32OiW
B1G1ER4CWg4dT1kgxqGg+Hj8ibDUiMFRMXU6rR6D3I63vKS21KHwfYCDdb0l8KTr
+2MY0wZ+Nz5Ya0tgrBE1T1VxmM/ccjEAjErgipb9K5fKaiNJMU0HCysrlBB5KTNX
0e7K93GLTAc+qkCyD0guXHN9q/YtnNzNjA+oQLH4F+v7dQaUzUZbxMcULQ+qG/vG
flaoFUexxxT0yL7gAlLS1bMqRjGLkwX8WT+e3SkIK2VxIqDbxeIa9X6C4pf+p9/d
BuizaE/58/WO/XQhOEyREcTZhwrNAt8Gf+z7EKM+ePEm6ygH/3B66zPu4d6BIJAA
R1lCcQZMbXmIXqEzi67JKX5O/UJMW7CW7X0mQwH0Kadv2UeHvRN+1uDNdXsGJ9vj
Ut8sIvpEFCRpXZpPWwbYkFk1+HOEKwmlb3Q1HioAQlLaCkricCwJquwLUCsv/9Jy
H6SUhKAW0m8rhQmJHI7Po4aIy3MmXOe8uajw4dvIgS7baz0g6jKgGDwwdaemsxCl
sJ6zz0C8xRD/xXaKMf8O484JZDkkAnmO2vr0d+r+yEpu3USd4Btf4rlu1jz3J5ct
jGAQNu+QMyfa85cBx5TD/l2UPiJntKrIFRhaj6ZFkDTIkLFkNgyAsiojvi0cONJP
AUZWdGUBrS9vMCgQAv1AdXfzcvJ1Uex0n+lJ+hfPcIm2NhKvoD9sMdPYR1O5Txfo
8vpfq6rvKV3heHVnBoOxhPt2iPeWEf/waOKIRePC891x8Te5ZtsKUa9Yl3yektX3
IfMzmJI38KkE9IUGQdNeS5ZwW07K9ScW3w1ckVAnkMSuDlRuGy35YGd3WppzWvUn
zLW1ZCTHC2/I318HTxYDUVwYBrho1Cri2fqhMu9VFX9PdSLSqMiGYDxGY/ktpqUT
/87CHCLh9MvOxB0HL31xTLP42Y9wlPsa47XfFRljwiRvoNiP+tLqW2ys1oDAelHP
5HJEy0jUGjJSa538OH6fa3O3qiWxyYqBr+99+3Hb7eXhSWiVBOuTtXaHm17ZAGs3
Whd/1HKqb2P0lkk9cNUTp84m5GIdDFkSUCdLtzX9Thd4Svsomtqg/sIXXaawsk//
qFWloZJIPz10nXTlLPcwAtIuXWTMpb/03U23LRqFEG2fOi5jYfQSVl6gvp+yWuZ2
BXaWXK7ghoUEAJU/N7k/IgGSXM5g9wOV6/NnyjWS1tTETiG2QGAHyXBb57c3kMHF
anEN6Nir4IsDuL7KWH1OBfPXQMhRn0RDftTxMNMHBkZii0DdutlLoOIdM9leUYig
ARTAlicbhKRTPLBNOqlrC+gCiFuvDjqvVbd6T3IgGP3Xe9RXoeKEvo/oiEV31yJF
l+Ln7tQVMivDusI0X6blT/o6LgElWI03i/a8LToi0vdRE1TFeZ/Q6ttIkdQIcZ8v
ptehFUGArPojRif0A161sgmnWsNavEuPxHPK3BFnExwiptqun/U6Hz0I1FBuREQj
BqdQ5ojZb0mP39E+Cbx4RGC0y5gR6MVuPtaTNA2FYed2+KvgDQxgm4d1hRhBbDxG
zwpvp7n2IN51RaG5JEHYGltcM1AVhsdQC8RqJeAtR05meUlLMBazJki5WyBZDmrG
95KF76GNZHrMC9j9zSQgriP5ZHM+L4MHM9UaSBhwhyKWbnSCjxLN3/SKVDLU/f67
ovWGtRF+ZY/arqwxMM+EJE3CbBuaFyWxr+u5PlvpYBO3prBJMqaAISPOEOSgAXeQ
f8nEXR8Wfq5hvJRl+NRxKUyyBdICli8gdDWidNeBR2YP5ERbJg1lIXvwihz4XWCD
1KhffkRditlJDw3XR9dkhTuSyzqVd5iOk9C3hAQldOQ9GY1vh7ekRaySCcSS8wSp
Z0ZIVhHZiB8mVIre1t71NHvDaPLlPau6QtjSrCgF5yJKklBI3TBpqaAZzni8L31U
LtMT3tPShV0SgoZ1CnGxkwLI+POLrlKGVOpk2xlLAMIvh0UxgAy2z2FDbitqVDkL
GMUvegC0Q8PlZfqo/eM9uNK1Whv/z1N54juNMqc6gSZ/6OwstvT1CHhQQl3eu4II
8AlCfo6g+bTzrlMvMotQ3jRbCtaIS5S6AB4O6OhMOcdP55oKnwwn73sf47QLRTaY
WqubPgWZd5f2YW9a3TeEdV+jv5EMDqFutAUUFU9Tk0AlwP+NI+D9sJ3UUlL/Gebz
67g0iqsrAJEz56sJD+4SXI0ulw27AGsgFhElr+r3Vxz7eegi+UIDGMiE9hFRkSjY
7j9qzdEb5uV2PU7GZGCt1BcgtoJx6mt2OcwCnvyAhbz9LwepZVjHJQSlzi68iCsg
iz8Ya5f9JgCHR/Oax53bGJ9b4GsZVVqoLC93VcMblruyRDgVDPk858GZbjpVp6wS
VA4jYrc78XglYk2eoQcnPf0J3g27VADJRfpkBNwkct33L/JrOzp6SgIQQvjxi5Fx
5BVxoaUkHU6D1u3C6r7wtY7FjXIcvgslkI7JvM3WcChD51e/7HBQGrlqb9Akq9Xh
m7PdfPVAMuy87X6UunT8BLBjvmhvRAeeW9r21Be++Tbh1OqiVxAVF+14zRC3cbIe
3UrCKR3s34CAiW/mB8eIenKE2ZZcIV2H/79ZIhX+9LU0cuSqPa699Jiby3Ro1F+8
Pcmg0HquFnXHhw7MgL4HU9HKvnZNSe6PE5oNMZB/QgKVW/Fc5LiBcU3jSfsrD+Ae
a1aGVFB1Hst67kg2w+wPJrBZSqYe2oRpmQm1abn5lrdaNKnpOZsEYMOjgsEp6lpg
hVijEdBFoImzFtnIgyguaKSYhlc3+Lm4Mec8yVw4/d8o0jjw+eoaWNgRwVmO1xAN
cq3gqaitUtpYCXXWVQU38+eGDbfheGOuTjq7y2hK9HIX/PLdATItT+3rkWZYzYY5
s/fphp3jHY3pDfMZ3ib9ufixPtvkkPMhQJOsahSFTcDuvRsn42S02LpiRQ/Mfy8I
3Ed0vZUpOqVZ//FIsAtD1WhzkevU9qgufJXrLKpIZyvqVC4WU/qV2e3bdatYa4tZ
K2MR4VVTmEjo+BL+55DKjnzRyUsa6EzawfAsNtvwCpwP7VIVABusN0nrC+ZhxT2v
Pckvq2cYEm2bm3P7S1SoZhwvsCRInjmtIZTdthcd5S3bb2OrH7Xj7DEviF4sbcXM
SSvYb5bUG6NzMjTSDXiVzzqsg7e4v7sp3qVe7RMTBy91miKsbq9QlVszP0os/prE
Jb3z1jEobrYeCyfcJPYvXUXJPwZ3Fqi30nwjkYaBVKnPQWSNWhpJ49OMJx5DGa41
C8QEydQUTfNFM1AWzeGNAoddb7HPXTJjK4wiKHnR+rfUa+4sgIHzERYrpzlFAC7q
35PDqvtmukZh9JWd/Imvpw0YZVfx1fvc2t2945WeSiRmNqpK52IIP4vowSgU1zy/
ZzGB3c3vvYAeJISWdREZkC7CNtvY1wsxc3fOC5PtDl0Owf8yulKTmafAopayRfHL
5ASWvK8DaQjqFE5+SnO9xt4ksdUICFBKITpblBx+rw0nyYX+gusC1cTK7ckoGa/Q
XNhRSTK6I4hnfmQmO5gOBLwX2djwi0jMzK3bQoMGVa9fliyJDcXQOsHqpl1s5Ref
JtNsTQth7tfvtJvvYQI0Qw+gwQzmwWC8o/q2tgCLsf8bJ84mX376kX5vUWt6300R
40QYDY2+45RpsL+HprqGGGSOIJvr93oze/iDNpqTUw5suPdNZoqZNvVXClwVoHdY
bvwIFsNTY3d0ovoPZNURNgi3QmdlMJUfuaVGROM2Sdpz3TJhRH+ZRLQh1tOapmm2
X7UGjPk99q3zmpKbrM0rreYZWppQK5ZR04xMBCcgaZxWfFq4zBBPeTK+9P/OO8K+
YDopwX6JTo3E6bbDk1SD1ciBR0bxERwzaJbPq5n92oWCHaCim+YAa6IQ/Zdzm25N
fTyAkxfTSqr3bXtqMDHTIwkMoQm2kq4py3cCnEpyycjjwO2DCBlg6Y9QfIHYqmQi
2KRRpyGU9q3Q+6pHbbuIVyi63yiRqxgKZkT69Ki2+uPJGq4uEeKXcPGgjGUxewA5
yhJwVt9/wGeIMAoqQxGGYoISIPvukrpYOiNk99mNMfx+ZiLZxOKxglwO/o28gMhp
/cshElV3elSKAXt+uvo92XjYmMxviWiRHB3JFiSboY2L+KY3AMOnJKIozFcnWGeg
bVzk3mC5QNVhW8h9LMm7L4MZx7xc/huWt7s6qKgK6ZUHudO3jIMnc4iX0NkJGLGB
77id+sP+X22w5XTygLtx+r2t7CfEsTsK0VJEaewVFTNLWtv03nlvnuhn8tEaQacf
Wh4ofTBjzLhIuXGlEHsQeKoxwmUC6hjBK0aRRpiMc2XZpIvGb0ZkKJ2k9LUOktSv
VPhIdVu73FNYHqg1R6IF4BTe/7NNSSvwW1ifSIGrmqcHyLeq3oHV93tF68CTNoq0
lF8sSXXi/5Ws9BUImMyNoqReVg2ozNQkHF9Lcm5stFc0XLKVCLJjDv+S/ynauXpZ
MYZ+0wARzKCBPQKk9GLmfY7eijyJA2SdN+3siHqf9DGG5HsqTH+hH9CkvuqAfbqr
xY4Gojq7YekXT30QHFLHxvg/xYWk9PIyGd+0LXZ68VAjrw7BLlu+Eg7pt7i1r5Mo
OXzUmZ391pjk3VzT1zJgXuB7A30yvEY4nT06vaViXy66H2u92ku84TJqJEkRO4Hz
NSoqRRDEHM0aGfccfUZWef1UYKu7ix3EAVWI6/MTjNniJ3N+UIgE8xGl+qtKE2nc
AGkjYYSeTAiaQzZ8mx6EX5VKmMOfxo0/UlSlJrCvbPPh5iFAR37ElkZvDy5baAie
XC4oNukJRSJsmU92EwYg8yozt38zTzz3nKB8sV/p+KUM+uGisGR3eHX/45KUgmQi
G55R/ylVwYeL7xZY0dBDW5vhI5n4epY5yr+FTenkaTVLweZtb1dhYwVQ3PwQtEU0
qx8+nMTH8TrvxiVHDC5Gd2loa65tgBG/2wD8WizThWUvr8b9kGqus4Zno1Zs57u8
O6zLcC6Ka18td2/CyavgbbLFj/Ti7fX5MBfiB0QHX1RkVtqQpag1zIeQ15eGSipt
5JJMcITOL+KsrLGveTqa08eTC7Fho+CYv1R+aSpfR2uy2l2JF+daukur+is4RQTc
/NdYmfVM5zlBRPitLdefJmitoCNqzTiEKBEKS3jjhThr75ZD5ADhllFknzV+VM3u
T+gylDDZ/LcEToUEhvEnR9ZUZ52wnUlUGkvND7F9cgHT0v7AhznjXxtjWB9cIrh0
h9j4/S4TsAbHfz14cjylOAoXU/+37IPln8wHzrxP2Duh1Pads0+ztfQlrEz4QdoZ
qO8DMtfydQsH1JJnkALz4TJSO8wAowESxfBWPYfYcpR7Tfmy5JpmXoulFj7g5nm/
ITYl6TcEtEhUx78CN3YO1UML58EhLc6R46yE2ARovUA9hd3Laef6odoYM12rl1UA
95MtjTmiAtNAIcNOn3msyAqDvbhFxSO2GkF/3kIbJ4CwJVPfeSqOn5/AUEEVMFBQ
OzjbiSNhEFQaAk5lSkZzFJTlfNVY2jG0HOrb77SwxiRxWXPeIbYYVpawojoXQKha
vPLQdxGsiu02M7Q4hJNPkW4z+BQ+DHjRF/NKhbZiOveURAmeOgo15REYEQnCu4R5
yzCdLIRkj03bIbqdwQwbgevler2jCYPpW9MrGWkxN9vynO/7AS3jV499KG9xPeaU
LD4cxENdjvEt0sDZSShaIJ5t6uhoUYLVAcxIWXS8UizKyPhjET3HU7IAqJrux+4e
nfXjjKrJeVGVyxW600I1ovhVdwmwYkkErH+nQZa6nQnK4OIU/KLUtqtBlyIpM18u
fzkZgWpftAM/Km8sYvVGETfECJ5vG2ll+QiZgen85VEmsCTGm0zSKaclJCFWOjex
D80rdZ0lulpoLTOAcGHxyGqsnN/1z/69F6WbtC2g8q+9QK1Toun8M47Wvcgy5opk
yNbqm0PM2Dw50eTiKoN2oy2xs//8jKkxkuWfXISJXwiISFZ35oc3YOj1KzYlKQsy
T4cs1sEXSQ02ERZJWireeQHvk7YOLpwgmZyzWVMjxwkiDvKz/m6b8m8mo3zbdt85
BLq3GMho3tGmVSC4Js+ew8sr230HfM+ckteFYolh2PU+mQ4eQ/sj4oi5qqBVE5U6
OVG99FnhcHAM8E9Lqb+Y7g8lDK/lATsw/GGmgmpGCzhAewDIXp63g1qL/6G/3y4q
5zKw/T5qrt+8KbrcNsbyBvWkYU3eg6j8oduxF3o7vUhQL8wf+Yj3+kR06Uina3t+
mEo4gA06Scg6wnuyE8Otssjr9RWdni+3vOgC4/8W1Y8Yu8Cs0o29RO/QT1vuH6I1
eYrNFMZ7x/G9knkmSTVQ8ENo7x3bJ3H2gKnSlVsnTP63UhRT+94ltlm54UcuQugA
y7HRa7nFJlhdaJoOf2deEEBt+43z0FskEcJCNmGCFH+wA3zJIWzioK8896QEUGYv
fdVPNxrJL0HrgOt3UkOlVZOfExksNyj2yCiS2sl1c/9oJwa1Tf7dZOxYaNJQv29O
NrZLbn0e9WQzmKVzy3t5JE+yCMm5/sFuUuRxMt3YefUJVVktx3Zd6MVB/4PkVVI6
zAJM2nDATqKphyspAS1X25IkAW71fvyYW2SLJzxzlY7ufWz6kJHwwPhbuy/4qHou
6GG/35i13Fm4q5q1OvlATFhkpkOXLvJiH4Mz8X11l1UXh7vis1fzYAnXyv+vktBE
gmJli559ZIbLXYmERn7cCWxG0YU7h/+VpxdbJGjEoJR4pT4QOr8pNMATMJVqaDXC
Vi6odHU3MOEUqgTEwjaUnXoGU3L8OVXYYg/TZ19ScQrn34GuGcdrzlfKJKpWN0p7
Ih7mpuJA9dRtson71kzAdIQlYIZmFlxaVNEIIpR/bjdf2ILzi0qrg5fDihhxOpZO
I4M1P1LRJIJ2Qg097S58fraUUnoyfrYmD4oFWCWoCZOAVPRzoGHZEFTSfLZSAE3o
FuKBqjvP7i3vKZGblL+4dc7au4GMQ2Qa4zrx+2SaxJR4KmTlvL3rtsC7ulDYe7yA
j8HXi4lruiYVX6qNRRU7JtlMFvRUlpIICZTddf9sHtKnyLj39h9L5RpOujv1hOjF
Bn73hrDd2ZPVRHowFBiCysTTaF56/qOxU/y5n/qj0nla1YkZBlJ/ik0TyL879/o3
3NNdhTrzge7bdUCwDJ7VAoOgr/otTrNYPVngqkDA19Rs2T4kUkkUhiMXILiUa93U
+J0slVw+4x5gJnuDQEwksUWX1Vhu2eUgU/mEbcBZ69X2c5GAFK2NKGO3AAzuEm/p
rPRvHlFe0rvwpHHjLwl1w9cEA2p4J4M+A0Hiq8W40kCxp0i0oB8kiQnAQqL3N3hP
tAod2m0PG8bb/gFmiWiIpXwzqmGkhFR8BhVEIXAoLbPS5/1EnKOmiTVVBF+9xsQS
vjoR9fR3fejOAn0V5ppvFo3cYN/ahq1c8Y2GrMuq+lNK3YCQj6BT0fR2J9ONhtYg
HWvJ4ZdO+MlZOJc37P3E/Usv40lWnRKXAt5VAY1L2SxWXy5XIdiOcE5gL8ssB/mq
pG9jDRomuS87+dqAhpxA472P6V4isGA48td9Z2NVloawMgE1Yl22sTFaTd1/uxGG
stmSeRNggRO685pBCU1meSXsuN/mU2JlppQvohqmKGKc1e4c2iwJM1EnqMnAhxFq
HHg4W0JJSbPZqe0FWT9AK0nxkYPk/VARoCENUU9mXWLo1/pcvuLiPTCYhUDiBXCv
uHIFYahvX7X0F8NR4/8f51VdWIBQH5bLWMp1UOjia3B+WSCubh5SqhgvX1KMEJjN
V+k0sPN7esZHi1KqGcZJ7pf9O7bryfEIvajuEDdo0QxNdZaB+JI4qD81q6wOZr//
OEhd4Y5jZbspPitcVXDWDIcDly1pJMmlZHbnTzbeK1HjSC8kazzhk0t+Zxbf61h1
AbA2ZIFSnB35GOpwB0IX8B1khTOnEMcX+gSQ5vyiQXm9UdY67wXsT0VrK04vzliX
uF68wDls8vuURPFbbQT0dTHDaHAdGoDubpyv1W+uKGAEXIf7s7MaWl57up6vbhU+
wFjM4Q7lsYXAioOsTKlToKE9cQ0XZNu3D39CXYFEKx0w0xg1cLvmrZTVDGaGB4a4
UjLsRUltEf9jvMREKgCLmQfxaCH5jLMCvap1tM9zpOE5B8f0kn1j22Y53QsoS45A
gyNywePO4SZ6XQdDYNNOD8V7r9IibPhejo+wLsSM6rPqEaM91Idluwl/ZExFq1JI
5onUkvEin6mArBXnmZDUdpT70nOeZlMVf2KHVx7t2IFvlNSJ0F9YU0Daa6ar/+y+
gWd+cU3kBcHsTajGLTgxjk5BdAOJG9jVEIAf2yIAsuh9T2wgVKmtiU64rD7mq0Xd
+qjNbetWpt51olZ08wxZuz8F5EZuKsZxDqe8/Yf4SNAJkvvOpyLK4EZk6dz3NZQ4
x7qBaz7zUtR8V4sQDJ2tHIXfTvrPjMm5gnAhHDnfSvyYwSafbrxl5IllqMiQlOTQ
q4BYaR3ECfDJ/XCY82VoJUBJ2rLWs8vdV0WVaDK55q+2YMTtFK1tFOTSXogNk9+v
WZwhhPViznP7d/ZZMGBWdBdFms2BvFWbEuUSliii3b7+NDFmLlfmcXw8d3oASt7d
G4dVsL7RMwHsiNgqlHuiQ/2vvBl46WIuCmVcd/R2S9/mT6qZr/LAvu3KEAlRnMfr
uvzuk4ZAygwZJvF2i+qydJR9hbLHCPhZQ9DLvk3o6KdT82RCrM5tydYWlmupKMGM
KyUJySzSCfmw3t06ctd3GsrYkSjwjiMjoB1yabzgIajHNzIQc9wkK3XF81EDlJ3F
NQZaVLYeYDJA39cIBXknh6oHpBhOtQr5vu1qBqbBVxJ5gOkAFHH+0jADTvnXkVzG
VC1lD58bZgLXqGVdaxLbuM11elZYZPX+hUVPGlzqQDgve+FYOxNeGYklLvt0eNKm
slpCDTN+oDrgW8sYBK69YkL8/G2d7+i+GejQafhL7Gk/BDjCr2++WY2occr78U4I
2wE0qVeLk7eNzuSyRvimCi+sJlYQWF2ZYQHdfDDyBa1tyUvEZjj1gmqzDxKa4G1j
pMy4dZWK2/oOrcBcvlg0hx6le7yg3CTpV2TftzN8KYI5oobNEFs7jcSWAVJ/wS53
rjn7O0HYO+VT7T5cqf7c5OZs5kSt6UHgeolncubMCKP0+IaMa0D6t3xwq5R5XihJ
4VnOziG8yL4YdKyxTCL4gIeMaDBxgrmS7RYHT6bFM78vqlLL0EduIECAY0V1bcbW
FyDsbGk9x4JQjdvbAEbYXzoTWeI79H8l4u4k5MbyekduY6XDzhhFTe7WoZ90HB6P
xj3Fevnk+bFeVE0mR3RFbTrWO7s4x2uGCfHTZY+QzBQ9I4zXSYbcqCwksmjUWgC4
Sg78+qdC/gEPNg4uxx1aJ6Xf5fAqXQYZ5UVzFdLkWWIUSGLJp8KzsYJbZwHPxQ0n
BhYEo5EutSCJW0/BP/4u9ZOlNDd+CTTEx5M9DmxkbD6zfrUAW3mTZFRye/Ursqpn
9sZ38cqskUZ5HVvZUG080mVar0ZzkNncpfXc5++IM8Gwke7XDoeMdtGgeHIlSe6o
jfM3gkTv2GnrxK8+uenehQ0OxheL4j1zZWxjE/AxKiBf2Q2bZW19+b7jYlGcG7/8
qTTAxMX3QQWPJ7wtOZvoruBa5hKWxxSygghAQO058ZA6oVYStCPV9xOpFG8/uPZT
KPURmjsz10bozX/6ojIwSHMKXTjl1yd8Vw8NqNQB0QppfJRA2iaIpUuoSmBEV9/P
XzI1WmObzLDZcMxc3L/00O5vBieAEqsJIg4p7fVdKcPsclvo7VMmkYiDXUBkTZ+P
zwmKDAGpY6drisZAX27uwee27XF62SlbiPJNqL1udY5T5zy+UxgaDbPcTYKwbkfJ
R512hecw7E/L2uDvsoRqI5/yVmSTGV4AW2O3S69VZGP96kV9uND+/WYAYo+0ucNr
VNX8b/OGYBgtpB8p8twGssx7jqcrHr0IwNo7EA9Jonv5vbnJHHYtbokgzgS4q93e
XOPUz9htEaFNDLCofvc/5f/y3NXVFa35fyAObnJSagAw2kA9Ls9KqZNMdP7P3/I7
Nxjj89oMwfqF7nwt2gjGlHMCmJpBN30KE5y1gUZ3W0RpgvSdI3bk7bt36fMt4Y5m
vrmO0P6TsG3+nLMfqmMFoWNuVO7w6IHFvbGcbOTRChHxMorKshZPWOrulZbXy/H2
ukOI+0vM1BoAEWtt9TpF/v+cPClUrpyqreXbKt1AQK88Q/34Kgx4jVm5dop9sQD/
zhkUjIVZuGieO53IpdsbyKlYpFDW0ZqelUmf+C88opJDQiEfqTwprDI5QWDbFXVe
7bcyZwVBf0ukb/gvgqgw4RaQfmbhwq8uvZel8UssZw3PTjz6DEoYHR4Du+idGS0p
kFVU6gB8cvzqLHEXDMbioX3DdAQUxLCLTMD6nnIv/jzE/iJthdNy8+Y2occV2/18
jOr7/xEXVrCztWhHV/zgztKVqfh1RPEO08wKrY05wZAG5Z4BQMYdpb/eiX73XU5Q
eBCkgwoGwcdGkapSgCNDr0pb4J8l+TemlfI4rytbrFKZ4jJNnrS4an7D8LrLFUur
BLd8EXQw4mXSZJ06OWN8DW7+Ab1gFToSgGds6alypdgTkuHx6MksinU2GXuF7SeZ
s8waSBMgI/rSlr78gsDvaczEf8Q6gpiq9UB3/Jq66m73kHBXbQNMnNPzmb7+xwCD
JFCai4xqvNWjCTx5FPnGLXtw3HpdFo+Jto3XMb+IYH9i9iL0XrTUJCDhWH25pRrH
S7/jgF09nuxdmgqvYQO5mpM7sqnZPzOGCGdorYYwi5Uz2pGn6oJdYF3hmwoRTQM8
J8BTZ/mwOZE7l7h3kc3Q8rmCcfvIn9pr2DXkaaI5dN2R8ZDZ++pnh+eAWFNey4d5
pxfMX0T2gK8paPiNQfUcijZyG4pm41/+NXKrjK91eSvk1SuhtZz0EM4HtVZTpOeb
uqVY65ZP62TefUCzO7zbrK7MIKRbVTBBv28bjIA5OtoBpRdGYFNtjXZrefo9SFQC
TDbovO+J1s33A3l5iWEqbZ2ObRYNe2dPqWbM+4DUICr+/ETVIDWdXHNS8RuSIA0e
Lu+zEv4Gy3p1Jm0a6nODhuySnP7rQINTsQDq2FN7BdCbDFuTQkza+Dv8RH1LErTT
aX6nQj/G9Zy8zz/vEgYwePX1yvUc7X4rkniNN/IcayvUWzR0hs4IZJGSoxcEeKaZ
Uu/3Q9vLhAKCWG96Tykp+4sSKl6CrudFTnzymG6ucbebg16YoKDbxTet/hSLCGff
stBEz7WDVbMbW/n+s6EsRANShBaIru/wca8+kzy0HrP/zfCo8SstTi3jF4Kuud6L
XRWfH7jjjd0ZvdQT7IN4FHIA/ItzsRx55BheNkYpjuHwAVKMqbk7leH5MtvWpJkR
aU3DwVbK9UG36i6p+UXHOpzd0KxmhvGxgHBURFODlS0HrUOMeLBYwZkNDmmujC9f
leCLfv23R8gcCZgxFNq+5enUgsWprAbgA4+T9ZX444hkIYfnLZdVjC2nDGNx984X
O3mUX+vnuoNEmmIUkVo4xugRHKHsuT68/hCkA+oMW17+2d3SjUVyJVyhf6DysrRU
6v5PKxI0OMY/hfmMhbvajsASKGkYEeL8JvOtsyZQ/h7/V3l7DoSUs4nqhFL0XOj0
ID+7okNiXNt3l7w8zkMePL+j5HJ9nI/Guj0yRUSzMTXo8LxcNOM5ICXPqlPAUo9w
ajG+dJ+rM0vR+QU5gqkg1S81P/Be17M3j69abmQF73mkLafXwFoUyKqrg+J61MfE
L616hhVoXCouk3sabZZkmx8K43xIeoD6HDJGb+UOED4NVaLRLGoi1azZ4f+OjdW7
Ej98xBPR6B2KbxqV0jj4Rxso8KESDdcv8Pv7YJ42SsMNkVZyBmiiHrCL3bqnHN4W
POa9owAC9W8YkVUJexr0lglnHo65uTHQ5+IpDwWX81+5+pCCl1I6/+FzHQfBbW+y
77ArBqfdTVKop9QNfT8aU+QQfLfpx/a3AugUNnQzskERuQCK5gwThJUHU/07M22f
zvsGOOU6ryIeBOS1JxegDsGMQP+gTgdRf71Er9RiJnYIJLFsKdSXbKWexANOMkhi
bB4Ri94/W8yFktgffxrZMZZxFMivaApLu5erAvSN9ax0jCrxTRsKGRcPFh+qjLQw
PGWLcfhNpniPn/hok9dPRbhrrzovPGLwP3gyDE6oH5rrzZSZYME/LmZD19l8UMjV
nCaxhg+dN7t1j/m3GXS4CL7jJgGqo3lnt6EKEqvO4kIEP+ng1e8+XhGRfrWj3t8H
4qxD2mhDehG90ZBb+dEE0bqtAVz7YOwyIopE2TJgz2df50Z9GnlfAQ0Rq2xdWvVn
VfaGgx7EF6SAgFaeE4S+LVjBKIFu4qka/zjy9kPcWlaADZx7SsBTL/Il7CqpDD2S
vIz1E28Yp8nFb6rJ2TbcSw33y3Sob071+1bBxWJA16yzO7Fxw4czVzgCFmAGj5lr
3kT2niT8JSwDvGA4mYexwbUfcKGJZ12Qsl9CdYFPAjes5vcgcWbNSgUu4/mdoa9+
NwiaJ095jC+tqsAyBQEyRhrfLg+6RflErdiky9yrmFUsVU2Lqr70z1S47n2wfC8i
uJafAXWnh7SV8poOpULhB5MSAbXbDgCv4aBxlYVtWbgXMJKoSYfz7PTFmypmcvME
Iw6ASctCC1XXsFw4Q1KGjVbgYQ4mw0oTv2ABT5qYs3QLANBCoVC5pkWCI4GT+OcT
WZ+gYdcCwrwJ4VmT384PyzXHxmIcKU6IPcC4999htgEmtP5kvGaq+R+FGLBKGA0K
m6a9OfgYmR+ks67vb2S5u+QJrYJRpeNt43paAokP4gC4lYUndVyWV3VXYEEk5Fol
UX1uagCncfn9A8xIH9bo8B29OML77Go1Hc5LKq0A55SYsqCJgx8Sf1mi70KBx3pU
GMxde4mNk6SXEKn5ILSRBwaLWv9kdKVbmydbGfjf+yU0Kdtwv9w46gofnMsqC8kL
3u+bjorBlQ25udmr3T9AzujaaOGTcMwJM3gxI8c/I+Scj7wFgK1ceMjrx39LG8KQ
f1QKhodqeT8TobZ+Wog8153tX1kjfyyl3q7TCQJL2dZM410EaMxJNXYN4Amd/c71
mCceGY0f0Q6kM8UBVAQTFof+bOoBOOnTxKCb6uc0WD5wv1ZgjSCnLy19esHcv4J9
9aKFL2shGegmTOAiqgmnmLH5srs6fseh7ZPzVfI+aEi2MRFVXgNASfl/L3u2PbcC
LFXxhhBVgngv9t3qPezQsWgqaPqIq/IPSDRffklqLGctHWahTI/6e/y9PwY5lFxM
zRFJNHR18hP29Kx2pQCFZN33oq4kRZOnOW/VmFrwxPIevHGgHjy5gbEzWNnlTYFb
M7nawVrr/g3C82IP0dP+jiqDUYn/sgfPGArGx/Do6fk81sUPGt9WI66JA6NsSa2M
95UCJCssIjc4iq8e33LQbdaVo1/PyPKAiF93VKHhKRt9PXzqF11qVYMhvVZNVP05
xop6u32yqXI1MsscoCYyhoXe1ji0c7wyuUtTyTg41yHKy6gH6+deCAxmzigLdPdb
/Dvf2nwiEwMSIOXF6dnnBHMReQfeX6k7IPO8zEuAL/+vSyIc+0XncrGgalcS2N7r
XUI5cAr4sYthzkmhlYiduaQklO1C4v/nWDA1C88QEIc23u1K2zeZ8zi9Yuw1RAMo
OHh2fR+zT+Co4tW4NUh7XBrgJPXWzdF6eO0v0IvmY69GWGdVGAxle4x17Z3IjIdm
SVeiUG2sZH8s7fkM8wWigMFbEm4yOZ/IkRZAZgsBsyc/6UQMu4DcBq7ZmgTiTAxY
+BP5+Ol6Q1NQ9BnCqbb/76fDysjfUnxx3mxMoQELZiPZYu+3O//quXF/RvN5QQBq
PIC78AlmqQrc8vasbEOQ9X/saRGlTrceovc44CGAPN+I+Q6ivUGsnfYDQymUqYLC
KY6oj7be8C7SXx9jD0UqWf5mwnx1CNizbtpKZkp951HGBQYXHo/kNsrEsRnAh5Hu
4hVw4IQ39WiZ0ctpGY/VQKpYhaTRyeBkL+1d7bG6FdFCMA0K5pGqtYLjCr9ORGU+
gmg3Mi5kRMxtB69oDCLQA6qyvobrgjxDTvj+rVOdEuiqvErRcsomda8TVDTwDAfK
xK5jxCKDxt4iBHa2EN2/GrEDUY4H6xV2iGpX5DPgV4o28oKcfn7YBmak/la5UI/P
fumyodBaAS5ztSznGsqRV+2C0B3+NHlMi+kfR8KJ1cy2RiX8WYZfWkYTb/5zYuOA
MJBrddSnYk5viVbef4up5QmcEqxsAOsy/+jkZ9aNN0cBrs0KlDpG9amgwhM4k2en
rU6DDMqybacGbIW6N9F1checyOCIkSFPcG026H8BhCLCRwgK8b7NCVYq6CsruVvv
Dpp2bVG2bpwGCDTYcc8giFqTFdnZ0Aq8qNbUUhIsyJRld5KeYPZciVz6Mt5ETLKZ
6UV0KlnLKaItGfbl5jVKyCFrp9bqwinBmBKhnc3nvmjSPsyPyxp2DfVe0aGihCCz
nNoWf9tolR/XDL5Tyal1muR2Gt/QP5ZTlXn0ylBBqf3puPtaXaMdYyz4bIsFvTIy
7dxUGwR4wp23vKjgMvOg6jEvwrmVlte9nhjUMEg5l2E2ZI//d7Xh09/iI5TL6RAA
p3R54lgpCxP8EIuMmkJfyd4iPWmsT26rQOVasaslh/1D8UKjuJOadLmOriWymviD
1Vb6nv9zJm+JWyDHXT1P+rag8Myr3Odb0JGQD9YPJVh4f1V3rZqIAX+Mhqs6oGlc
8qiRQsRphOtrwW2ZaJ7DzwqBc8tlBleEVIleUZ6MDJOoGLjWvtWO7jiOt24OsBoI
Qq9GMAVasmVxY6Wlhe/N1AdzhVFSBBEbB5rNWUoeqlaSYzWL4N7LAUtUh80HwEGK
4HcjK5pBGvHXEp3HcmmtwDomq8c5K7gpaLmrVVrWZnOMQ9QreQyeKEKgt2KrLvg0
iMkxdhZqlHK1KGkjWtgC4a3t2V9DxV9KOR1gBDEKfS+jHHfNbKfeYUirgjLz5RRj
eM6yz+yEjRt2OZlimkHABOwlZYWWq9DIxByU0tCXlKT1CGR55a+R7zNGUaY8ajyl
U1G40CJXb7Cc8f7biNyl305dWpqmnhwYJDOua6GpF+ZYC4xEL4mR1hwZZH0OycWG
GKgE0/XqcBdGw4U2jAIORGXu5E/vbbkDLcYhSk9IE122X0WrKm3FL8Y/EjykAN4P
7Qo+FjcaoOzWPCjkSluaC+RcM2UVPGUso77fSuNc8Zbw8o6Ufn1vH3HhKauTWyzH
hMLR89QPQMP5o02QLfqH84zA5zMGzMwremxePgXPB0ipmcfnIlMdzstatkGkcyjb
vEfT0lggVJeXU1mO+93ScFRjV1Ogn3iftj6z69zpWzWiLXWEb4RyGUIVLErsZdfp
05VLEFtXTUL5t5t0mX/NDhR6mb1B5CK0Nrh6lKpBSLamKLdm5tel4EY226a/81uv
PKP8/TohpYwonwrFOzTMjLRol3zMa/xsqRoJax8xOjokz1mfa9jpJm+VCFQHZxz3
lN/hk9B3QeiaiDqyjRyOLaupxAL7lrbp0lMLhH5wzDUGJ9yHVr5pzA1bvg/TxU2K
hjuduiW/Z2r4OxhccQzzyOmNF6TRsDHGVFju/u5pFFCC+qoVLADd9HoPugvhbu8d
eildxReVtvILankDozldwAPRayMkVTf+Y/yPSPX4NhqMcffDaUHcsWbjsg9k5pdX
hZGxMHdHwYQ1UK7xvwvRbOjWZ8WLErYmCp04JRJru/Hco0s/W4Sxgzj19zfARwNI
8lWm0nOwE40LXmNt8xTMcK8uCZi+Cf79Xo9VdFYjoh0wX3uGdhb2TIN6PMyMNcim
mtPz9QfAEA4xC+OUGkKN2th+x7Vfk+QXO48P7PpcfvTXXtD3DEbMCmMJ+Se8IdSV
JUEpvM02dbMZ1/+nr8DG9pAr1Tnd22EZWws0k1+JdblC7gZNnr305NPQlcMkuejE
dHazLOQcFlBTOgeDajtbEin7WQz8TvpfYIXy+DgqY4/6UwxIo2Tcl+Gm5PZk8Vik
FWas4lZfkNbzLNpNwYvpwKVdDif/lOAbxk4+p83tY4Z3dKl9cHLJCegWHUsaOWYE
G+Q+vdSUiX23DImrJdxKy4ooDd0vT+C9r9Y2rHc8FQzlnCDTncxNPS+2DbMppswm
8w2h7F0UnDWMnU8siyKKDtM6PZX+7VcoyyHD9uCaIvfLESzsLd8IVICCud9975T9
d9dOpft8w2Ns05jcOfMTNytq2hzLO+uc9JbDqRufGt5h0/WQstSLDYIPvepewonR
IH5tsbxxaSng9bLePz0ixpnsvbz9oyZ/GR8uWUUHO8l1x+O8VG/ACm6/B1MXY+/4
dLb3F7k/Knz7VbRN/3/UIz+0m0aFfXkSBt6FuEBgVDo+GvJb6Oh3pMULnxDG98ID
VnTHv+JEblCIsEHsJWDowTqDXpJNGB1AGg37apWH0tSRwYzEWkcxZbAr/bOEx1TH
tmWf+JUTUOwLEUsx1px/Sm2Lbn4n3CsekKopfVThK7VOEjpE9h8KMk3ZO19S0aOw
lCgbt4dJhCgMsKcw2xs5fw6Dy4ik0W1JkISIH5qCunqv6755Xefeqd0S9sMDRETY
NshGKU1A3hLfCmDBN7djnDLjsAVfwlnWhrf34ZHBP4cZjRJIxGO3vcT88NwkW+d6
ss87SVGSbfIHi30hyHZyFII4vGozooJXPiQ+4h9frT/L38Y1RnJdu+77J6PJxvjJ
M1paRV4dytoLHxX6srl4hKYs6eh3+aeN8Gar8mxRYz0=
`protect end_protected
